module QuireToPosit256_16_0(
  input          clock,
  input          reset,
  input          io_inValid,
  input  [313:0] io_quireIn,
  output [15:0]  io_positOut,
  output         io_outValid
);
  wire [312:0] _T; // @[QuireToPosit.scala 47:43]
  wire  _T_1; // @[QuireToPosit.scala 47:47]
  wire  tailIsZero; // @[QuireToPosit.scala 47:27]
  wire  _T_2; // @[QuireToPosit.scala 49:45]
  wire  outRawFloat_isNaR; // @[QuireToPosit.scala 49:49]
  wire  _T_5; // @[QuireToPosit.scala 50:31]
  wire  outRawFloat_isZero; // @[QuireToPosit.scala 50:51]
  wire [312:0] _T_8; // @[QuireToPosit.scala 58:41]
  wire [312:0] _T_9; // @[QuireToPosit.scala 58:68]
  wire [312:0] quireXOR; // @[QuireToPosit.scala 58:56]
  wire [255:0] _T_10; // @[LZD.scala 43:32]
  wire [127:0] _T_11; // @[LZD.scala 43:32]
  wire [63:0] _T_12; // @[LZD.scala 43:32]
  wire [31:0] _T_13; // @[LZD.scala 43:32]
  wire [15:0] _T_14; // @[LZD.scala 43:32]
  wire [7:0] _T_15; // @[LZD.scala 43:32]
  wire [3:0] _T_16; // @[LZD.scala 43:32]
  wire [1:0] _T_17; // @[LZD.scala 43:32]
  wire  _T_18; // @[LZD.scala 39:14]
  wire  _T_19; // @[LZD.scala 39:21]
  wire  _T_20; // @[LZD.scala 39:30]
  wire  _T_21; // @[LZD.scala 39:27]
  wire  _T_22; // @[LZD.scala 39:25]
  wire [1:0] _T_23; // @[Cat.scala 29:58]
  wire [1:0] _T_24; // @[LZD.scala 44:32]
  wire  _T_25; // @[LZD.scala 39:14]
  wire  _T_26; // @[LZD.scala 39:21]
  wire  _T_27; // @[LZD.scala 39:30]
  wire  _T_28; // @[LZD.scala 39:27]
  wire  _T_29; // @[LZD.scala 39:25]
  wire [1:0] _T_30; // @[Cat.scala 29:58]
  wire  _T_31; // @[Shift.scala 12:21]
  wire  _T_32; // @[Shift.scala 12:21]
  wire  _T_33; // @[LZD.scala 49:16]
  wire  _T_34; // @[LZD.scala 49:27]
  wire  _T_35; // @[LZD.scala 49:25]
  wire  _T_36; // @[LZD.scala 49:47]
  wire  _T_37; // @[LZD.scala 49:59]
  wire  _T_38; // @[LZD.scala 49:35]
  wire [2:0] _T_40; // @[Cat.scala 29:58]
  wire [3:0] _T_41; // @[LZD.scala 44:32]
  wire [1:0] _T_42; // @[LZD.scala 43:32]
  wire  _T_43; // @[LZD.scala 39:14]
  wire  _T_44; // @[LZD.scala 39:21]
  wire  _T_45; // @[LZD.scala 39:30]
  wire  _T_46; // @[LZD.scala 39:27]
  wire  _T_47; // @[LZD.scala 39:25]
  wire [1:0] _T_48; // @[Cat.scala 29:58]
  wire [1:0] _T_49; // @[LZD.scala 44:32]
  wire  _T_50; // @[LZD.scala 39:14]
  wire  _T_51; // @[LZD.scala 39:21]
  wire  _T_52; // @[LZD.scala 39:30]
  wire  _T_53; // @[LZD.scala 39:27]
  wire  _T_54; // @[LZD.scala 39:25]
  wire [1:0] _T_55; // @[Cat.scala 29:58]
  wire  _T_56; // @[Shift.scala 12:21]
  wire  _T_57; // @[Shift.scala 12:21]
  wire  _T_58; // @[LZD.scala 49:16]
  wire  _T_59; // @[LZD.scala 49:27]
  wire  _T_60; // @[LZD.scala 49:25]
  wire  _T_61; // @[LZD.scala 49:47]
  wire  _T_62; // @[LZD.scala 49:59]
  wire  _T_63; // @[LZD.scala 49:35]
  wire [2:0] _T_65; // @[Cat.scala 29:58]
  wire  _T_66; // @[Shift.scala 12:21]
  wire  _T_67; // @[Shift.scala 12:21]
  wire  _T_68; // @[LZD.scala 49:16]
  wire  _T_69; // @[LZD.scala 49:27]
  wire  _T_70; // @[LZD.scala 49:25]
  wire [1:0] _T_71; // @[LZD.scala 49:47]
  wire [1:0] _T_72; // @[LZD.scala 49:59]
  wire [1:0] _T_73; // @[LZD.scala 49:35]
  wire [3:0] _T_75; // @[Cat.scala 29:58]
  wire [7:0] _T_76; // @[LZD.scala 44:32]
  wire [3:0] _T_77; // @[LZD.scala 43:32]
  wire [1:0] _T_78; // @[LZD.scala 43:32]
  wire  _T_79; // @[LZD.scala 39:14]
  wire  _T_80; // @[LZD.scala 39:21]
  wire  _T_81; // @[LZD.scala 39:30]
  wire  _T_82; // @[LZD.scala 39:27]
  wire  _T_83; // @[LZD.scala 39:25]
  wire [1:0] _T_84; // @[Cat.scala 29:58]
  wire [1:0] _T_85; // @[LZD.scala 44:32]
  wire  _T_86; // @[LZD.scala 39:14]
  wire  _T_87; // @[LZD.scala 39:21]
  wire  _T_88; // @[LZD.scala 39:30]
  wire  _T_89; // @[LZD.scala 39:27]
  wire  _T_90; // @[LZD.scala 39:25]
  wire [1:0] _T_91; // @[Cat.scala 29:58]
  wire  _T_92; // @[Shift.scala 12:21]
  wire  _T_93; // @[Shift.scala 12:21]
  wire  _T_94; // @[LZD.scala 49:16]
  wire  _T_95; // @[LZD.scala 49:27]
  wire  _T_96; // @[LZD.scala 49:25]
  wire  _T_97; // @[LZD.scala 49:47]
  wire  _T_98; // @[LZD.scala 49:59]
  wire  _T_99; // @[LZD.scala 49:35]
  wire [2:0] _T_101; // @[Cat.scala 29:58]
  wire [3:0] _T_102; // @[LZD.scala 44:32]
  wire [1:0] _T_103; // @[LZD.scala 43:32]
  wire  _T_104; // @[LZD.scala 39:14]
  wire  _T_105; // @[LZD.scala 39:21]
  wire  _T_106; // @[LZD.scala 39:30]
  wire  _T_107; // @[LZD.scala 39:27]
  wire  _T_108; // @[LZD.scala 39:25]
  wire [1:0] _T_109; // @[Cat.scala 29:58]
  wire [1:0] _T_110; // @[LZD.scala 44:32]
  wire  _T_111; // @[LZD.scala 39:14]
  wire  _T_112; // @[LZD.scala 39:21]
  wire  _T_113; // @[LZD.scala 39:30]
  wire  _T_114; // @[LZD.scala 39:27]
  wire  _T_115; // @[LZD.scala 39:25]
  wire [1:0] _T_116; // @[Cat.scala 29:58]
  wire  _T_117; // @[Shift.scala 12:21]
  wire  _T_118; // @[Shift.scala 12:21]
  wire  _T_119; // @[LZD.scala 49:16]
  wire  _T_120; // @[LZD.scala 49:27]
  wire  _T_121; // @[LZD.scala 49:25]
  wire  _T_122; // @[LZD.scala 49:47]
  wire  _T_123; // @[LZD.scala 49:59]
  wire  _T_124; // @[LZD.scala 49:35]
  wire [2:0] _T_126; // @[Cat.scala 29:58]
  wire  _T_127; // @[Shift.scala 12:21]
  wire  _T_128; // @[Shift.scala 12:21]
  wire  _T_129; // @[LZD.scala 49:16]
  wire  _T_130; // @[LZD.scala 49:27]
  wire  _T_131; // @[LZD.scala 49:25]
  wire [1:0] _T_132; // @[LZD.scala 49:47]
  wire [1:0] _T_133; // @[LZD.scala 49:59]
  wire [1:0] _T_134; // @[LZD.scala 49:35]
  wire [3:0] _T_136; // @[Cat.scala 29:58]
  wire  _T_137; // @[Shift.scala 12:21]
  wire  _T_138; // @[Shift.scala 12:21]
  wire  _T_139; // @[LZD.scala 49:16]
  wire  _T_140; // @[LZD.scala 49:27]
  wire  _T_141; // @[LZD.scala 49:25]
  wire [2:0] _T_142; // @[LZD.scala 49:47]
  wire [2:0] _T_143; // @[LZD.scala 49:59]
  wire [2:0] _T_144; // @[LZD.scala 49:35]
  wire [4:0] _T_146; // @[Cat.scala 29:58]
  wire [15:0] _T_147; // @[LZD.scala 44:32]
  wire [7:0] _T_148; // @[LZD.scala 43:32]
  wire [3:0] _T_149; // @[LZD.scala 43:32]
  wire [1:0] _T_150; // @[LZD.scala 43:32]
  wire  _T_151; // @[LZD.scala 39:14]
  wire  _T_152; // @[LZD.scala 39:21]
  wire  _T_153; // @[LZD.scala 39:30]
  wire  _T_154; // @[LZD.scala 39:27]
  wire  _T_155; // @[LZD.scala 39:25]
  wire [1:0] _T_156; // @[Cat.scala 29:58]
  wire [1:0] _T_157; // @[LZD.scala 44:32]
  wire  _T_158; // @[LZD.scala 39:14]
  wire  _T_159; // @[LZD.scala 39:21]
  wire  _T_160; // @[LZD.scala 39:30]
  wire  _T_161; // @[LZD.scala 39:27]
  wire  _T_162; // @[LZD.scala 39:25]
  wire [1:0] _T_163; // @[Cat.scala 29:58]
  wire  _T_164; // @[Shift.scala 12:21]
  wire  _T_165; // @[Shift.scala 12:21]
  wire  _T_166; // @[LZD.scala 49:16]
  wire  _T_167; // @[LZD.scala 49:27]
  wire  _T_168; // @[LZD.scala 49:25]
  wire  _T_169; // @[LZD.scala 49:47]
  wire  _T_170; // @[LZD.scala 49:59]
  wire  _T_171; // @[LZD.scala 49:35]
  wire [2:0] _T_173; // @[Cat.scala 29:58]
  wire [3:0] _T_174; // @[LZD.scala 44:32]
  wire [1:0] _T_175; // @[LZD.scala 43:32]
  wire  _T_176; // @[LZD.scala 39:14]
  wire  _T_177; // @[LZD.scala 39:21]
  wire  _T_178; // @[LZD.scala 39:30]
  wire  _T_179; // @[LZD.scala 39:27]
  wire  _T_180; // @[LZD.scala 39:25]
  wire [1:0] _T_181; // @[Cat.scala 29:58]
  wire [1:0] _T_182; // @[LZD.scala 44:32]
  wire  _T_183; // @[LZD.scala 39:14]
  wire  _T_184; // @[LZD.scala 39:21]
  wire  _T_185; // @[LZD.scala 39:30]
  wire  _T_186; // @[LZD.scala 39:27]
  wire  _T_187; // @[LZD.scala 39:25]
  wire [1:0] _T_188; // @[Cat.scala 29:58]
  wire  _T_189; // @[Shift.scala 12:21]
  wire  _T_190; // @[Shift.scala 12:21]
  wire  _T_191; // @[LZD.scala 49:16]
  wire  _T_192; // @[LZD.scala 49:27]
  wire  _T_193; // @[LZD.scala 49:25]
  wire  _T_194; // @[LZD.scala 49:47]
  wire  _T_195; // @[LZD.scala 49:59]
  wire  _T_196; // @[LZD.scala 49:35]
  wire [2:0] _T_198; // @[Cat.scala 29:58]
  wire  _T_199; // @[Shift.scala 12:21]
  wire  _T_200; // @[Shift.scala 12:21]
  wire  _T_201; // @[LZD.scala 49:16]
  wire  _T_202; // @[LZD.scala 49:27]
  wire  _T_203; // @[LZD.scala 49:25]
  wire [1:0] _T_204; // @[LZD.scala 49:47]
  wire [1:0] _T_205; // @[LZD.scala 49:59]
  wire [1:0] _T_206; // @[LZD.scala 49:35]
  wire [3:0] _T_208; // @[Cat.scala 29:58]
  wire [7:0] _T_209; // @[LZD.scala 44:32]
  wire [3:0] _T_210; // @[LZD.scala 43:32]
  wire [1:0] _T_211; // @[LZD.scala 43:32]
  wire  _T_212; // @[LZD.scala 39:14]
  wire  _T_213; // @[LZD.scala 39:21]
  wire  _T_214; // @[LZD.scala 39:30]
  wire  _T_215; // @[LZD.scala 39:27]
  wire  _T_216; // @[LZD.scala 39:25]
  wire [1:0] _T_217; // @[Cat.scala 29:58]
  wire [1:0] _T_218; // @[LZD.scala 44:32]
  wire  _T_219; // @[LZD.scala 39:14]
  wire  _T_220; // @[LZD.scala 39:21]
  wire  _T_221; // @[LZD.scala 39:30]
  wire  _T_222; // @[LZD.scala 39:27]
  wire  _T_223; // @[LZD.scala 39:25]
  wire [1:0] _T_224; // @[Cat.scala 29:58]
  wire  _T_225; // @[Shift.scala 12:21]
  wire  _T_226; // @[Shift.scala 12:21]
  wire  _T_227; // @[LZD.scala 49:16]
  wire  _T_228; // @[LZD.scala 49:27]
  wire  _T_229; // @[LZD.scala 49:25]
  wire  _T_230; // @[LZD.scala 49:47]
  wire  _T_231; // @[LZD.scala 49:59]
  wire  _T_232; // @[LZD.scala 49:35]
  wire [2:0] _T_234; // @[Cat.scala 29:58]
  wire [3:0] _T_235; // @[LZD.scala 44:32]
  wire [1:0] _T_236; // @[LZD.scala 43:32]
  wire  _T_237; // @[LZD.scala 39:14]
  wire  _T_238; // @[LZD.scala 39:21]
  wire  _T_239; // @[LZD.scala 39:30]
  wire  _T_240; // @[LZD.scala 39:27]
  wire  _T_241; // @[LZD.scala 39:25]
  wire [1:0] _T_242; // @[Cat.scala 29:58]
  wire [1:0] _T_243; // @[LZD.scala 44:32]
  wire  _T_244; // @[LZD.scala 39:14]
  wire  _T_245; // @[LZD.scala 39:21]
  wire  _T_246; // @[LZD.scala 39:30]
  wire  _T_247; // @[LZD.scala 39:27]
  wire  _T_248; // @[LZD.scala 39:25]
  wire [1:0] _T_249; // @[Cat.scala 29:58]
  wire  _T_250; // @[Shift.scala 12:21]
  wire  _T_251; // @[Shift.scala 12:21]
  wire  _T_252; // @[LZD.scala 49:16]
  wire  _T_253; // @[LZD.scala 49:27]
  wire  _T_254; // @[LZD.scala 49:25]
  wire  _T_255; // @[LZD.scala 49:47]
  wire  _T_256; // @[LZD.scala 49:59]
  wire  _T_257; // @[LZD.scala 49:35]
  wire [2:0] _T_259; // @[Cat.scala 29:58]
  wire  _T_260; // @[Shift.scala 12:21]
  wire  _T_261; // @[Shift.scala 12:21]
  wire  _T_262; // @[LZD.scala 49:16]
  wire  _T_263; // @[LZD.scala 49:27]
  wire  _T_264; // @[LZD.scala 49:25]
  wire [1:0] _T_265; // @[LZD.scala 49:47]
  wire [1:0] _T_266; // @[LZD.scala 49:59]
  wire [1:0] _T_267; // @[LZD.scala 49:35]
  wire [3:0] _T_269; // @[Cat.scala 29:58]
  wire  _T_270; // @[Shift.scala 12:21]
  wire  _T_271; // @[Shift.scala 12:21]
  wire  _T_272; // @[LZD.scala 49:16]
  wire  _T_273; // @[LZD.scala 49:27]
  wire  _T_274; // @[LZD.scala 49:25]
  wire [2:0] _T_275; // @[LZD.scala 49:47]
  wire [2:0] _T_276; // @[LZD.scala 49:59]
  wire [2:0] _T_277; // @[LZD.scala 49:35]
  wire [4:0] _T_279; // @[Cat.scala 29:58]
  wire  _T_280; // @[Shift.scala 12:21]
  wire  _T_281; // @[Shift.scala 12:21]
  wire  _T_282; // @[LZD.scala 49:16]
  wire  _T_283; // @[LZD.scala 49:27]
  wire  _T_284; // @[LZD.scala 49:25]
  wire [3:0] _T_285; // @[LZD.scala 49:47]
  wire [3:0] _T_286; // @[LZD.scala 49:59]
  wire [3:0] _T_287; // @[LZD.scala 49:35]
  wire [5:0] _T_289; // @[Cat.scala 29:58]
  wire [31:0] _T_290; // @[LZD.scala 44:32]
  wire [15:0] _T_291; // @[LZD.scala 43:32]
  wire [7:0] _T_292; // @[LZD.scala 43:32]
  wire [3:0] _T_293; // @[LZD.scala 43:32]
  wire [1:0] _T_294; // @[LZD.scala 43:32]
  wire  _T_295; // @[LZD.scala 39:14]
  wire  _T_296; // @[LZD.scala 39:21]
  wire  _T_297; // @[LZD.scala 39:30]
  wire  _T_298; // @[LZD.scala 39:27]
  wire  _T_299; // @[LZD.scala 39:25]
  wire [1:0] _T_300; // @[Cat.scala 29:58]
  wire [1:0] _T_301; // @[LZD.scala 44:32]
  wire  _T_302; // @[LZD.scala 39:14]
  wire  _T_303; // @[LZD.scala 39:21]
  wire  _T_304; // @[LZD.scala 39:30]
  wire  _T_305; // @[LZD.scala 39:27]
  wire  _T_306; // @[LZD.scala 39:25]
  wire [1:0] _T_307; // @[Cat.scala 29:58]
  wire  _T_308; // @[Shift.scala 12:21]
  wire  _T_309; // @[Shift.scala 12:21]
  wire  _T_310; // @[LZD.scala 49:16]
  wire  _T_311; // @[LZD.scala 49:27]
  wire  _T_312; // @[LZD.scala 49:25]
  wire  _T_313; // @[LZD.scala 49:47]
  wire  _T_314; // @[LZD.scala 49:59]
  wire  _T_315; // @[LZD.scala 49:35]
  wire [2:0] _T_317; // @[Cat.scala 29:58]
  wire [3:0] _T_318; // @[LZD.scala 44:32]
  wire [1:0] _T_319; // @[LZD.scala 43:32]
  wire  _T_320; // @[LZD.scala 39:14]
  wire  _T_321; // @[LZD.scala 39:21]
  wire  _T_322; // @[LZD.scala 39:30]
  wire  _T_323; // @[LZD.scala 39:27]
  wire  _T_324; // @[LZD.scala 39:25]
  wire [1:0] _T_325; // @[Cat.scala 29:58]
  wire [1:0] _T_326; // @[LZD.scala 44:32]
  wire  _T_327; // @[LZD.scala 39:14]
  wire  _T_328; // @[LZD.scala 39:21]
  wire  _T_329; // @[LZD.scala 39:30]
  wire  _T_330; // @[LZD.scala 39:27]
  wire  _T_331; // @[LZD.scala 39:25]
  wire [1:0] _T_332; // @[Cat.scala 29:58]
  wire  _T_333; // @[Shift.scala 12:21]
  wire  _T_334; // @[Shift.scala 12:21]
  wire  _T_335; // @[LZD.scala 49:16]
  wire  _T_336; // @[LZD.scala 49:27]
  wire  _T_337; // @[LZD.scala 49:25]
  wire  _T_338; // @[LZD.scala 49:47]
  wire  _T_339; // @[LZD.scala 49:59]
  wire  _T_340; // @[LZD.scala 49:35]
  wire [2:0] _T_342; // @[Cat.scala 29:58]
  wire  _T_343; // @[Shift.scala 12:21]
  wire  _T_344; // @[Shift.scala 12:21]
  wire  _T_345; // @[LZD.scala 49:16]
  wire  _T_346; // @[LZD.scala 49:27]
  wire  _T_347; // @[LZD.scala 49:25]
  wire [1:0] _T_348; // @[LZD.scala 49:47]
  wire [1:0] _T_349; // @[LZD.scala 49:59]
  wire [1:0] _T_350; // @[LZD.scala 49:35]
  wire [3:0] _T_352; // @[Cat.scala 29:58]
  wire [7:0] _T_353; // @[LZD.scala 44:32]
  wire [3:0] _T_354; // @[LZD.scala 43:32]
  wire [1:0] _T_355; // @[LZD.scala 43:32]
  wire  _T_356; // @[LZD.scala 39:14]
  wire  _T_357; // @[LZD.scala 39:21]
  wire  _T_358; // @[LZD.scala 39:30]
  wire  _T_359; // @[LZD.scala 39:27]
  wire  _T_360; // @[LZD.scala 39:25]
  wire [1:0] _T_361; // @[Cat.scala 29:58]
  wire [1:0] _T_362; // @[LZD.scala 44:32]
  wire  _T_363; // @[LZD.scala 39:14]
  wire  _T_364; // @[LZD.scala 39:21]
  wire  _T_365; // @[LZD.scala 39:30]
  wire  _T_366; // @[LZD.scala 39:27]
  wire  _T_367; // @[LZD.scala 39:25]
  wire [1:0] _T_368; // @[Cat.scala 29:58]
  wire  _T_369; // @[Shift.scala 12:21]
  wire  _T_370; // @[Shift.scala 12:21]
  wire  _T_371; // @[LZD.scala 49:16]
  wire  _T_372; // @[LZD.scala 49:27]
  wire  _T_373; // @[LZD.scala 49:25]
  wire  _T_374; // @[LZD.scala 49:47]
  wire  _T_375; // @[LZD.scala 49:59]
  wire  _T_376; // @[LZD.scala 49:35]
  wire [2:0] _T_378; // @[Cat.scala 29:58]
  wire [3:0] _T_379; // @[LZD.scala 44:32]
  wire [1:0] _T_380; // @[LZD.scala 43:32]
  wire  _T_381; // @[LZD.scala 39:14]
  wire  _T_382; // @[LZD.scala 39:21]
  wire  _T_383; // @[LZD.scala 39:30]
  wire  _T_384; // @[LZD.scala 39:27]
  wire  _T_385; // @[LZD.scala 39:25]
  wire [1:0] _T_386; // @[Cat.scala 29:58]
  wire [1:0] _T_387; // @[LZD.scala 44:32]
  wire  _T_388; // @[LZD.scala 39:14]
  wire  _T_389; // @[LZD.scala 39:21]
  wire  _T_390; // @[LZD.scala 39:30]
  wire  _T_391; // @[LZD.scala 39:27]
  wire  _T_392; // @[LZD.scala 39:25]
  wire [1:0] _T_393; // @[Cat.scala 29:58]
  wire  _T_394; // @[Shift.scala 12:21]
  wire  _T_395; // @[Shift.scala 12:21]
  wire  _T_396; // @[LZD.scala 49:16]
  wire  _T_397; // @[LZD.scala 49:27]
  wire  _T_398; // @[LZD.scala 49:25]
  wire  _T_399; // @[LZD.scala 49:47]
  wire  _T_400; // @[LZD.scala 49:59]
  wire  _T_401; // @[LZD.scala 49:35]
  wire [2:0] _T_403; // @[Cat.scala 29:58]
  wire  _T_404; // @[Shift.scala 12:21]
  wire  _T_405; // @[Shift.scala 12:21]
  wire  _T_406; // @[LZD.scala 49:16]
  wire  _T_407; // @[LZD.scala 49:27]
  wire  _T_408; // @[LZD.scala 49:25]
  wire [1:0] _T_409; // @[LZD.scala 49:47]
  wire [1:0] _T_410; // @[LZD.scala 49:59]
  wire [1:0] _T_411; // @[LZD.scala 49:35]
  wire [3:0] _T_413; // @[Cat.scala 29:58]
  wire  _T_414; // @[Shift.scala 12:21]
  wire  _T_415; // @[Shift.scala 12:21]
  wire  _T_416; // @[LZD.scala 49:16]
  wire  _T_417; // @[LZD.scala 49:27]
  wire  _T_418; // @[LZD.scala 49:25]
  wire [2:0] _T_419; // @[LZD.scala 49:47]
  wire [2:0] _T_420; // @[LZD.scala 49:59]
  wire [2:0] _T_421; // @[LZD.scala 49:35]
  wire [4:0] _T_423; // @[Cat.scala 29:58]
  wire [15:0] _T_424; // @[LZD.scala 44:32]
  wire [7:0] _T_425; // @[LZD.scala 43:32]
  wire [3:0] _T_426; // @[LZD.scala 43:32]
  wire [1:0] _T_427; // @[LZD.scala 43:32]
  wire  _T_428; // @[LZD.scala 39:14]
  wire  _T_429; // @[LZD.scala 39:21]
  wire  _T_430; // @[LZD.scala 39:30]
  wire  _T_431; // @[LZD.scala 39:27]
  wire  _T_432; // @[LZD.scala 39:25]
  wire [1:0] _T_433; // @[Cat.scala 29:58]
  wire [1:0] _T_434; // @[LZD.scala 44:32]
  wire  _T_435; // @[LZD.scala 39:14]
  wire  _T_436; // @[LZD.scala 39:21]
  wire  _T_437; // @[LZD.scala 39:30]
  wire  _T_438; // @[LZD.scala 39:27]
  wire  _T_439; // @[LZD.scala 39:25]
  wire [1:0] _T_440; // @[Cat.scala 29:58]
  wire  _T_441; // @[Shift.scala 12:21]
  wire  _T_442; // @[Shift.scala 12:21]
  wire  _T_443; // @[LZD.scala 49:16]
  wire  _T_444; // @[LZD.scala 49:27]
  wire  _T_445; // @[LZD.scala 49:25]
  wire  _T_446; // @[LZD.scala 49:47]
  wire  _T_447; // @[LZD.scala 49:59]
  wire  _T_448; // @[LZD.scala 49:35]
  wire [2:0] _T_450; // @[Cat.scala 29:58]
  wire [3:0] _T_451; // @[LZD.scala 44:32]
  wire [1:0] _T_452; // @[LZD.scala 43:32]
  wire  _T_453; // @[LZD.scala 39:14]
  wire  _T_454; // @[LZD.scala 39:21]
  wire  _T_455; // @[LZD.scala 39:30]
  wire  _T_456; // @[LZD.scala 39:27]
  wire  _T_457; // @[LZD.scala 39:25]
  wire [1:0] _T_458; // @[Cat.scala 29:58]
  wire [1:0] _T_459; // @[LZD.scala 44:32]
  wire  _T_460; // @[LZD.scala 39:14]
  wire  _T_461; // @[LZD.scala 39:21]
  wire  _T_462; // @[LZD.scala 39:30]
  wire  _T_463; // @[LZD.scala 39:27]
  wire  _T_464; // @[LZD.scala 39:25]
  wire [1:0] _T_465; // @[Cat.scala 29:58]
  wire  _T_466; // @[Shift.scala 12:21]
  wire  _T_467; // @[Shift.scala 12:21]
  wire  _T_468; // @[LZD.scala 49:16]
  wire  _T_469; // @[LZD.scala 49:27]
  wire  _T_470; // @[LZD.scala 49:25]
  wire  _T_471; // @[LZD.scala 49:47]
  wire  _T_472; // @[LZD.scala 49:59]
  wire  _T_473; // @[LZD.scala 49:35]
  wire [2:0] _T_475; // @[Cat.scala 29:58]
  wire  _T_476; // @[Shift.scala 12:21]
  wire  _T_477; // @[Shift.scala 12:21]
  wire  _T_478; // @[LZD.scala 49:16]
  wire  _T_479; // @[LZD.scala 49:27]
  wire  _T_480; // @[LZD.scala 49:25]
  wire [1:0] _T_481; // @[LZD.scala 49:47]
  wire [1:0] _T_482; // @[LZD.scala 49:59]
  wire [1:0] _T_483; // @[LZD.scala 49:35]
  wire [3:0] _T_485; // @[Cat.scala 29:58]
  wire [7:0] _T_486; // @[LZD.scala 44:32]
  wire [3:0] _T_487; // @[LZD.scala 43:32]
  wire [1:0] _T_488; // @[LZD.scala 43:32]
  wire  _T_489; // @[LZD.scala 39:14]
  wire  _T_490; // @[LZD.scala 39:21]
  wire  _T_491; // @[LZD.scala 39:30]
  wire  _T_492; // @[LZD.scala 39:27]
  wire  _T_493; // @[LZD.scala 39:25]
  wire [1:0] _T_494; // @[Cat.scala 29:58]
  wire [1:0] _T_495; // @[LZD.scala 44:32]
  wire  _T_496; // @[LZD.scala 39:14]
  wire  _T_497; // @[LZD.scala 39:21]
  wire  _T_498; // @[LZD.scala 39:30]
  wire  _T_499; // @[LZD.scala 39:27]
  wire  _T_500; // @[LZD.scala 39:25]
  wire [1:0] _T_501; // @[Cat.scala 29:58]
  wire  _T_502; // @[Shift.scala 12:21]
  wire  _T_503; // @[Shift.scala 12:21]
  wire  _T_504; // @[LZD.scala 49:16]
  wire  _T_505; // @[LZD.scala 49:27]
  wire  _T_506; // @[LZD.scala 49:25]
  wire  _T_507; // @[LZD.scala 49:47]
  wire  _T_508; // @[LZD.scala 49:59]
  wire  _T_509; // @[LZD.scala 49:35]
  wire [2:0] _T_511; // @[Cat.scala 29:58]
  wire [3:0] _T_512; // @[LZD.scala 44:32]
  wire [1:0] _T_513; // @[LZD.scala 43:32]
  wire  _T_514; // @[LZD.scala 39:14]
  wire  _T_515; // @[LZD.scala 39:21]
  wire  _T_516; // @[LZD.scala 39:30]
  wire  _T_517; // @[LZD.scala 39:27]
  wire  _T_518; // @[LZD.scala 39:25]
  wire [1:0] _T_519; // @[Cat.scala 29:58]
  wire [1:0] _T_520; // @[LZD.scala 44:32]
  wire  _T_521; // @[LZD.scala 39:14]
  wire  _T_522; // @[LZD.scala 39:21]
  wire  _T_523; // @[LZD.scala 39:30]
  wire  _T_524; // @[LZD.scala 39:27]
  wire  _T_525; // @[LZD.scala 39:25]
  wire [1:0] _T_526; // @[Cat.scala 29:58]
  wire  _T_527; // @[Shift.scala 12:21]
  wire  _T_528; // @[Shift.scala 12:21]
  wire  _T_529; // @[LZD.scala 49:16]
  wire  _T_530; // @[LZD.scala 49:27]
  wire  _T_531; // @[LZD.scala 49:25]
  wire  _T_532; // @[LZD.scala 49:47]
  wire  _T_533; // @[LZD.scala 49:59]
  wire  _T_534; // @[LZD.scala 49:35]
  wire [2:0] _T_536; // @[Cat.scala 29:58]
  wire  _T_537; // @[Shift.scala 12:21]
  wire  _T_538; // @[Shift.scala 12:21]
  wire  _T_539; // @[LZD.scala 49:16]
  wire  _T_540; // @[LZD.scala 49:27]
  wire  _T_541; // @[LZD.scala 49:25]
  wire [1:0] _T_542; // @[LZD.scala 49:47]
  wire [1:0] _T_543; // @[LZD.scala 49:59]
  wire [1:0] _T_544; // @[LZD.scala 49:35]
  wire [3:0] _T_546; // @[Cat.scala 29:58]
  wire  _T_547; // @[Shift.scala 12:21]
  wire  _T_548; // @[Shift.scala 12:21]
  wire  _T_549; // @[LZD.scala 49:16]
  wire  _T_550; // @[LZD.scala 49:27]
  wire  _T_551; // @[LZD.scala 49:25]
  wire [2:0] _T_552; // @[LZD.scala 49:47]
  wire [2:0] _T_553; // @[LZD.scala 49:59]
  wire [2:0] _T_554; // @[LZD.scala 49:35]
  wire [4:0] _T_556; // @[Cat.scala 29:58]
  wire  _T_557; // @[Shift.scala 12:21]
  wire  _T_558; // @[Shift.scala 12:21]
  wire  _T_559; // @[LZD.scala 49:16]
  wire  _T_560; // @[LZD.scala 49:27]
  wire  _T_561; // @[LZD.scala 49:25]
  wire [3:0] _T_562; // @[LZD.scala 49:47]
  wire [3:0] _T_563; // @[LZD.scala 49:59]
  wire [3:0] _T_564; // @[LZD.scala 49:35]
  wire [5:0] _T_566; // @[Cat.scala 29:58]
  wire  _T_567; // @[Shift.scala 12:21]
  wire  _T_568; // @[Shift.scala 12:21]
  wire  _T_569; // @[LZD.scala 49:16]
  wire  _T_570; // @[LZD.scala 49:27]
  wire  _T_571; // @[LZD.scala 49:25]
  wire [4:0] _T_572; // @[LZD.scala 49:47]
  wire [4:0] _T_573; // @[LZD.scala 49:59]
  wire [4:0] _T_574; // @[LZD.scala 49:35]
  wire [6:0] _T_576; // @[Cat.scala 29:58]
  wire [63:0] _T_577; // @[LZD.scala 44:32]
  wire [31:0] _T_578; // @[LZD.scala 43:32]
  wire [15:0] _T_579; // @[LZD.scala 43:32]
  wire [7:0] _T_580; // @[LZD.scala 43:32]
  wire [3:0] _T_581; // @[LZD.scala 43:32]
  wire [1:0] _T_582; // @[LZD.scala 43:32]
  wire  _T_583; // @[LZD.scala 39:14]
  wire  _T_584; // @[LZD.scala 39:21]
  wire  _T_585; // @[LZD.scala 39:30]
  wire  _T_586; // @[LZD.scala 39:27]
  wire  _T_587; // @[LZD.scala 39:25]
  wire [1:0] _T_588; // @[Cat.scala 29:58]
  wire [1:0] _T_589; // @[LZD.scala 44:32]
  wire  _T_590; // @[LZD.scala 39:14]
  wire  _T_591; // @[LZD.scala 39:21]
  wire  _T_592; // @[LZD.scala 39:30]
  wire  _T_593; // @[LZD.scala 39:27]
  wire  _T_594; // @[LZD.scala 39:25]
  wire [1:0] _T_595; // @[Cat.scala 29:58]
  wire  _T_596; // @[Shift.scala 12:21]
  wire  _T_597; // @[Shift.scala 12:21]
  wire  _T_598; // @[LZD.scala 49:16]
  wire  _T_599; // @[LZD.scala 49:27]
  wire  _T_600; // @[LZD.scala 49:25]
  wire  _T_601; // @[LZD.scala 49:47]
  wire  _T_602; // @[LZD.scala 49:59]
  wire  _T_603; // @[LZD.scala 49:35]
  wire [2:0] _T_605; // @[Cat.scala 29:58]
  wire [3:0] _T_606; // @[LZD.scala 44:32]
  wire [1:0] _T_607; // @[LZD.scala 43:32]
  wire  _T_608; // @[LZD.scala 39:14]
  wire  _T_609; // @[LZD.scala 39:21]
  wire  _T_610; // @[LZD.scala 39:30]
  wire  _T_611; // @[LZD.scala 39:27]
  wire  _T_612; // @[LZD.scala 39:25]
  wire [1:0] _T_613; // @[Cat.scala 29:58]
  wire [1:0] _T_614; // @[LZD.scala 44:32]
  wire  _T_615; // @[LZD.scala 39:14]
  wire  _T_616; // @[LZD.scala 39:21]
  wire  _T_617; // @[LZD.scala 39:30]
  wire  _T_618; // @[LZD.scala 39:27]
  wire  _T_619; // @[LZD.scala 39:25]
  wire [1:0] _T_620; // @[Cat.scala 29:58]
  wire  _T_621; // @[Shift.scala 12:21]
  wire  _T_622; // @[Shift.scala 12:21]
  wire  _T_623; // @[LZD.scala 49:16]
  wire  _T_624; // @[LZD.scala 49:27]
  wire  _T_625; // @[LZD.scala 49:25]
  wire  _T_626; // @[LZD.scala 49:47]
  wire  _T_627; // @[LZD.scala 49:59]
  wire  _T_628; // @[LZD.scala 49:35]
  wire [2:0] _T_630; // @[Cat.scala 29:58]
  wire  _T_631; // @[Shift.scala 12:21]
  wire  _T_632; // @[Shift.scala 12:21]
  wire  _T_633; // @[LZD.scala 49:16]
  wire  _T_634; // @[LZD.scala 49:27]
  wire  _T_635; // @[LZD.scala 49:25]
  wire [1:0] _T_636; // @[LZD.scala 49:47]
  wire [1:0] _T_637; // @[LZD.scala 49:59]
  wire [1:0] _T_638; // @[LZD.scala 49:35]
  wire [3:0] _T_640; // @[Cat.scala 29:58]
  wire [7:0] _T_641; // @[LZD.scala 44:32]
  wire [3:0] _T_642; // @[LZD.scala 43:32]
  wire [1:0] _T_643; // @[LZD.scala 43:32]
  wire  _T_644; // @[LZD.scala 39:14]
  wire  _T_645; // @[LZD.scala 39:21]
  wire  _T_646; // @[LZD.scala 39:30]
  wire  _T_647; // @[LZD.scala 39:27]
  wire  _T_648; // @[LZD.scala 39:25]
  wire [1:0] _T_649; // @[Cat.scala 29:58]
  wire [1:0] _T_650; // @[LZD.scala 44:32]
  wire  _T_651; // @[LZD.scala 39:14]
  wire  _T_652; // @[LZD.scala 39:21]
  wire  _T_653; // @[LZD.scala 39:30]
  wire  _T_654; // @[LZD.scala 39:27]
  wire  _T_655; // @[LZD.scala 39:25]
  wire [1:0] _T_656; // @[Cat.scala 29:58]
  wire  _T_657; // @[Shift.scala 12:21]
  wire  _T_658; // @[Shift.scala 12:21]
  wire  _T_659; // @[LZD.scala 49:16]
  wire  _T_660; // @[LZD.scala 49:27]
  wire  _T_661; // @[LZD.scala 49:25]
  wire  _T_662; // @[LZD.scala 49:47]
  wire  _T_663; // @[LZD.scala 49:59]
  wire  _T_664; // @[LZD.scala 49:35]
  wire [2:0] _T_666; // @[Cat.scala 29:58]
  wire [3:0] _T_667; // @[LZD.scala 44:32]
  wire [1:0] _T_668; // @[LZD.scala 43:32]
  wire  _T_669; // @[LZD.scala 39:14]
  wire  _T_670; // @[LZD.scala 39:21]
  wire  _T_671; // @[LZD.scala 39:30]
  wire  _T_672; // @[LZD.scala 39:27]
  wire  _T_673; // @[LZD.scala 39:25]
  wire [1:0] _T_674; // @[Cat.scala 29:58]
  wire [1:0] _T_675; // @[LZD.scala 44:32]
  wire  _T_676; // @[LZD.scala 39:14]
  wire  _T_677; // @[LZD.scala 39:21]
  wire  _T_678; // @[LZD.scala 39:30]
  wire  _T_679; // @[LZD.scala 39:27]
  wire  _T_680; // @[LZD.scala 39:25]
  wire [1:0] _T_681; // @[Cat.scala 29:58]
  wire  _T_682; // @[Shift.scala 12:21]
  wire  _T_683; // @[Shift.scala 12:21]
  wire  _T_684; // @[LZD.scala 49:16]
  wire  _T_685; // @[LZD.scala 49:27]
  wire  _T_686; // @[LZD.scala 49:25]
  wire  _T_687; // @[LZD.scala 49:47]
  wire  _T_688; // @[LZD.scala 49:59]
  wire  _T_689; // @[LZD.scala 49:35]
  wire [2:0] _T_691; // @[Cat.scala 29:58]
  wire  _T_692; // @[Shift.scala 12:21]
  wire  _T_693; // @[Shift.scala 12:21]
  wire  _T_694; // @[LZD.scala 49:16]
  wire  _T_695; // @[LZD.scala 49:27]
  wire  _T_696; // @[LZD.scala 49:25]
  wire [1:0] _T_697; // @[LZD.scala 49:47]
  wire [1:0] _T_698; // @[LZD.scala 49:59]
  wire [1:0] _T_699; // @[LZD.scala 49:35]
  wire [3:0] _T_701; // @[Cat.scala 29:58]
  wire  _T_702; // @[Shift.scala 12:21]
  wire  _T_703; // @[Shift.scala 12:21]
  wire  _T_704; // @[LZD.scala 49:16]
  wire  _T_705; // @[LZD.scala 49:27]
  wire  _T_706; // @[LZD.scala 49:25]
  wire [2:0] _T_707; // @[LZD.scala 49:47]
  wire [2:0] _T_708; // @[LZD.scala 49:59]
  wire [2:0] _T_709; // @[LZD.scala 49:35]
  wire [4:0] _T_711; // @[Cat.scala 29:58]
  wire [15:0] _T_712; // @[LZD.scala 44:32]
  wire [7:0] _T_713; // @[LZD.scala 43:32]
  wire [3:0] _T_714; // @[LZD.scala 43:32]
  wire [1:0] _T_715; // @[LZD.scala 43:32]
  wire  _T_716; // @[LZD.scala 39:14]
  wire  _T_717; // @[LZD.scala 39:21]
  wire  _T_718; // @[LZD.scala 39:30]
  wire  _T_719; // @[LZD.scala 39:27]
  wire  _T_720; // @[LZD.scala 39:25]
  wire [1:0] _T_721; // @[Cat.scala 29:58]
  wire [1:0] _T_722; // @[LZD.scala 44:32]
  wire  _T_723; // @[LZD.scala 39:14]
  wire  _T_724; // @[LZD.scala 39:21]
  wire  _T_725; // @[LZD.scala 39:30]
  wire  _T_726; // @[LZD.scala 39:27]
  wire  _T_727; // @[LZD.scala 39:25]
  wire [1:0] _T_728; // @[Cat.scala 29:58]
  wire  _T_729; // @[Shift.scala 12:21]
  wire  _T_730; // @[Shift.scala 12:21]
  wire  _T_731; // @[LZD.scala 49:16]
  wire  _T_732; // @[LZD.scala 49:27]
  wire  _T_733; // @[LZD.scala 49:25]
  wire  _T_734; // @[LZD.scala 49:47]
  wire  _T_735; // @[LZD.scala 49:59]
  wire  _T_736; // @[LZD.scala 49:35]
  wire [2:0] _T_738; // @[Cat.scala 29:58]
  wire [3:0] _T_739; // @[LZD.scala 44:32]
  wire [1:0] _T_740; // @[LZD.scala 43:32]
  wire  _T_741; // @[LZD.scala 39:14]
  wire  _T_742; // @[LZD.scala 39:21]
  wire  _T_743; // @[LZD.scala 39:30]
  wire  _T_744; // @[LZD.scala 39:27]
  wire  _T_745; // @[LZD.scala 39:25]
  wire [1:0] _T_746; // @[Cat.scala 29:58]
  wire [1:0] _T_747; // @[LZD.scala 44:32]
  wire  _T_748; // @[LZD.scala 39:14]
  wire  _T_749; // @[LZD.scala 39:21]
  wire  _T_750; // @[LZD.scala 39:30]
  wire  _T_751; // @[LZD.scala 39:27]
  wire  _T_752; // @[LZD.scala 39:25]
  wire [1:0] _T_753; // @[Cat.scala 29:58]
  wire  _T_754; // @[Shift.scala 12:21]
  wire  _T_755; // @[Shift.scala 12:21]
  wire  _T_756; // @[LZD.scala 49:16]
  wire  _T_757; // @[LZD.scala 49:27]
  wire  _T_758; // @[LZD.scala 49:25]
  wire  _T_759; // @[LZD.scala 49:47]
  wire  _T_760; // @[LZD.scala 49:59]
  wire  _T_761; // @[LZD.scala 49:35]
  wire [2:0] _T_763; // @[Cat.scala 29:58]
  wire  _T_764; // @[Shift.scala 12:21]
  wire  _T_765; // @[Shift.scala 12:21]
  wire  _T_766; // @[LZD.scala 49:16]
  wire  _T_767; // @[LZD.scala 49:27]
  wire  _T_768; // @[LZD.scala 49:25]
  wire [1:0] _T_769; // @[LZD.scala 49:47]
  wire [1:0] _T_770; // @[LZD.scala 49:59]
  wire [1:0] _T_771; // @[LZD.scala 49:35]
  wire [3:0] _T_773; // @[Cat.scala 29:58]
  wire [7:0] _T_774; // @[LZD.scala 44:32]
  wire [3:0] _T_775; // @[LZD.scala 43:32]
  wire [1:0] _T_776; // @[LZD.scala 43:32]
  wire  _T_777; // @[LZD.scala 39:14]
  wire  _T_778; // @[LZD.scala 39:21]
  wire  _T_779; // @[LZD.scala 39:30]
  wire  _T_780; // @[LZD.scala 39:27]
  wire  _T_781; // @[LZD.scala 39:25]
  wire [1:0] _T_782; // @[Cat.scala 29:58]
  wire [1:0] _T_783; // @[LZD.scala 44:32]
  wire  _T_784; // @[LZD.scala 39:14]
  wire  _T_785; // @[LZD.scala 39:21]
  wire  _T_786; // @[LZD.scala 39:30]
  wire  _T_787; // @[LZD.scala 39:27]
  wire  _T_788; // @[LZD.scala 39:25]
  wire [1:0] _T_789; // @[Cat.scala 29:58]
  wire  _T_790; // @[Shift.scala 12:21]
  wire  _T_791; // @[Shift.scala 12:21]
  wire  _T_792; // @[LZD.scala 49:16]
  wire  _T_793; // @[LZD.scala 49:27]
  wire  _T_794; // @[LZD.scala 49:25]
  wire  _T_795; // @[LZD.scala 49:47]
  wire  _T_796; // @[LZD.scala 49:59]
  wire  _T_797; // @[LZD.scala 49:35]
  wire [2:0] _T_799; // @[Cat.scala 29:58]
  wire [3:0] _T_800; // @[LZD.scala 44:32]
  wire [1:0] _T_801; // @[LZD.scala 43:32]
  wire  _T_802; // @[LZD.scala 39:14]
  wire  _T_803; // @[LZD.scala 39:21]
  wire  _T_804; // @[LZD.scala 39:30]
  wire  _T_805; // @[LZD.scala 39:27]
  wire  _T_806; // @[LZD.scala 39:25]
  wire [1:0] _T_807; // @[Cat.scala 29:58]
  wire [1:0] _T_808; // @[LZD.scala 44:32]
  wire  _T_809; // @[LZD.scala 39:14]
  wire  _T_810; // @[LZD.scala 39:21]
  wire  _T_811; // @[LZD.scala 39:30]
  wire  _T_812; // @[LZD.scala 39:27]
  wire  _T_813; // @[LZD.scala 39:25]
  wire [1:0] _T_814; // @[Cat.scala 29:58]
  wire  _T_815; // @[Shift.scala 12:21]
  wire  _T_816; // @[Shift.scala 12:21]
  wire  _T_817; // @[LZD.scala 49:16]
  wire  _T_818; // @[LZD.scala 49:27]
  wire  _T_819; // @[LZD.scala 49:25]
  wire  _T_820; // @[LZD.scala 49:47]
  wire  _T_821; // @[LZD.scala 49:59]
  wire  _T_822; // @[LZD.scala 49:35]
  wire [2:0] _T_824; // @[Cat.scala 29:58]
  wire  _T_825; // @[Shift.scala 12:21]
  wire  _T_826; // @[Shift.scala 12:21]
  wire  _T_827; // @[LZD.scala 49:16]
  wire  _T_828; // @[LZD.scala 49:27]
  wire  _T_829; // @[LZD.scala 49:25]
  wire [1:0] _T_830; // @[LZD.scala 49:47]
  wire [1:0] _T_831; // @[LZD.scala 49:59]
  wire [1:0] _T_832; // @[LZD.scala 49:35]
  wire [3:0] _T_834; // @[Cat.scala 29:58]
  wire  _T_835; // @[Shift.scala 12:21]
  wire  _T_836; // @[Shift.scala 12:21]
  wire  _T_837; // @[LZD.scala 49:16]
  wire  _T_838; // @[LZD.scala 49:27]
  wire  _T_839; // @[LZD.scala 49:25]
  wire [2:0] _T_840; // @[LZD.scala 49:47]
  wire [2:0] _T_841; // @[LZD.scala 49:59]
  wire [2:0] _T_842; // @[LZD.scala 49:35]
  wire [4:0] _T_844; // @[Cat.scala 29:58]
  wire  _T_845; // @[Shift.scala 12:21]
  wire  _T_846; // @[Shift.scala 12:21]
  wire  _T_847; // @[LZD.scala 49:16]
  wire  _T_848; // @[LZD.scala 49:27]
  wire  _T_849; // @[LZD.scala 49:25]
  wire [3:0] _T_850; // @[LZD.scala 49:47]
  wire [3:0] _T_851; // @[LZD.scala 49:59]
  wire [3:0] _T_852; // @[LZD.scala 49:35]
  wire [5:0] _T_854; // @[Cat.scala 29:58]
  wire [31:0] _T_855; // @[LZD.scala 44:32]
  wire [15:0] _T_856; // @[LZD.scala 43:32]
  wire [7:0] _T_857; // @[LZD.scala 43:32]
  wire [3:0] _T_858; // @[LZD.scala 43:32]
  wire [1:0] _T_859; // @[LZD.scala 43:32]
  wire  _T_860; // @[LZD.scala 39:14]
  wire  _T_861; // @[LZD.scala 39:21]
  wire  _T_862; // @[LZD.scala 39:30]
  wire  _T_863; // @[LZD.scala 39:27]
  wire  _T_864; // @[LZD.scala 39:25]
  wire [1:0] _T_865; // @[Cat.scala 29:58]
  wire [1:0] _T_866; // @[LZD.scala 44:32]
  wire  _T_867; // @[LZD.scala 39:14]
  wire  _T_868; // @[LZD.scala 39:21]
  wire  _T_869; // @[LZD.scala 39:30]
  wire  _T_870; // @[LZD.scala 39:27]
  wire  _T_871; // @[LZD.scala 39:25]
  wire [1:0] _T_872; // @[Cat.scala 29:58]
  wire  _T_873; // @[Shift.scala 12:21]
  wire  _T_874; // @[Shift.scala 12:21]
  wire  _T_875; // @[LZD.scala 49:16]
  wire  _T_876; // @[LZD.scala 49:27]
  wire  _T_877; // @[LZD.scala 49:25]
  wire  _T_878; // @[LZD.scala 49:47]
  wire  _T_879; // @[LZD.scala 49:59]
  wire  _T_880; // @[LZD.scala 49:35]
  wire [2:0] _T_882; // @[Cat.scala 29:58]
  wire [3:0] _T_883; // @[LZD.scala 44:32]
  wire [1:0] _T_884; // @[LZD.scala 43:32]
  wire  _T_885; // @[LZD.scala 39:14]
  wire  _T_886; // @[LZD.scala 39:21]
  wire  _T_887; // @[LZD.scala 39:30]
  wire  _T_888; // @[LZD.scala 39:27]
  wire  _T_889; // @[LZD.scala 39:25]
  wire [1:0] _T_890; // @[Cat.scala 29:58]
  wire [1:0] _T_891; // @[LZD.scala 44:32]
  wire  _T_892; // @[LZD.scala 39:14]
  wire  _T_893; // @[LZD.scala 39:21]
  wire  _T_894; // @[LZD.scala 39:30]
  wire  _T_895; // @[LZD.scala 39:27]
  wire  _T_896; // @[LZD.scala 39:25]
  wire [1:0] _T_897; // @[Cat.scala 29:58]
  wire  _T_898; // @[Shift.scala 12:21]
  wire  _T_899; // @[Shift.scala 12:21]
  wire  _T_900; // @[LZD.scala 49:16]
  wire  _T_901; // @[LZD.scala 49:27]
  wire  _T_902; // @[LZD.scala 49:25]
  wire  _T_903; // @[LZD.scala 49:47]
  wire  _T_904; // @[LZD.scala 49:59]
  wire  _T_905; // @[LZD.scala 49:35]
  wire [2:0] _T_907; // @[Cat.scala 29:58]
  wire  _T_908; // @[Shift.scala 12:21]
  wire  _T_909; // @[Shift.scala 12:21]
  wire  _T_910; // @[LZD.scala 49:16]
  wire  _T_911; // @[LZD.scala 49:27]
  wire  _T_912; // @[LZD.scala 49:25]
  wire [1:0] _T_913; // @[LZD.scala 49:47]
  wire [1:0] _T_914; // @[LZD.scala 49:59]
  wire [1:0] _T_915; // @[LZD.scala 49:35]
  wire [3:0] _T_917; // @[Cat.scala 29:58]
  wire [7:0] _T_918; // @[LZD.scala 44:32]
  wire [3:0] _T_919; // @[LZD.scala 43:32]
  wire [1:0] _T_920; // @[LZD.scala 43:32]
  wire  _T_921; // @[LZD.scala 39:14]
  wire  _T_922; // @[LZD.scala 39:21]
  wire  _T_923; // @[LZD.scala 39:30]
  wire  _T_924; // @[LZD.scala 39:27]
  wire  _T_925; // @[LZD.scala 39:25]
  wire [1:0] _T_926; // @[Cat.scala 29:58]
  wire [1:0] _T_927; // @[LZD.scala 44:32]
  wire  _T_928; // @[LZD.scala 39:14]
  wire  _T_929; // @[LZD.scala 39:21]
  wire  _T_930; // @[LZD.scala 39:30]
  wire  _T_931; // @[LZD.scala 39:27]
  wire  _T_932; // @[LZD.scala 39:25]
  wire [1:0] _T_933; // @[Cat.scala 29:58]
  wire  _T_934; // @[Shift.scala 12:21]
  wire  _T_935; // @[Shift.scala 12:21]
  wire  _T_936; // @[LZD.scala 49:16]
  wire  _T_937; // @[LZD.scala 49:27]
  wire  _T_938; // @[LZD.scala 49:25]
  wire  _T_939; // @[LZD.scala 49:47]
  wire  _T_940; // @[LZD.scala 49:59]
  wire  _T_941; // @[LZD.scala 49:35]
  wire [2:0] _T_943; // @[Cat.scala 29:58]
  wire [3:0] _T_944; // @[LZD.scala 44:32]
  wire [1:0] _T_945; // @[LZD.scala 43:32]
  wire  _T_946; // @[LZD.scala 39:14]
  wire  _T_947; // @[LZD.scala 39:21]
  wire  _T_948; // @[LZD.scala 39:30]
  wire  _T_949; // @[LZD.scala 39:27]
  wire  _T_950; // @[LZD.scala 39:25]
  wire [1:0] _T_951; // @[Cat.scala 29:58]
  wire [1:0] _T_952; // @[LZD.scala 44:32]
  wire  _T_953; // @[LZD.scala 39:14]
  wire  _T_954; // @[LZD.scala 39:21]
  wire  _T_955; // @[LZD.scala 39:30]
  wire  _T_956; // @[LZD.scala 39:27]
  wire  _T_957; // @[LZD.scala 39:25]
  wire [1:0] _T_958; // @[Cat.scala 29:58]
  wire  _T_959; // @[Shift.scala 12:21]
  wire  _T_960; // @[Shift.scala 12:21]
  wire  _T_961; // @[LZD.scala 49:16]
  wire  _T_962; // @[LZD.scala 49:27]
  wire  _T_963; // @[LZD.scala 49:25]
  wire  _T_964; // @[LZD.scala 49:47]
  wire  _T_965; // @[LZD.scala 49:59]
  wire  _T_966; // @[LZD.scala 49:35]
  wire [2:0] _T_968; // @[Cat.scala 29:58]
  wire  _T_969; // @[Shift.scala 12:21]
  wire  _T_970; // @[Shift.scala 12:21]
  wire  _T_971; // @[LZD.scala 49:16]
  wire  _T_972; // @[LZD.scala 49:27]
  wire  _T_973; // @[LZD.scala 49:25]
  wire [1:0] _T_974; // @[LZD.scala 49:47]
  wire [1:0] _T_975; // @[LZD.scala 49:59]
  wire [1:0] _T_976; // @[LZD.scala 49:35]
  wire [3:0] _T_978; // @[Cat.scala 29:58]
  wire  _T_979; // @[Shift.scala 12:21]
  wire  _T_980; // @[Shift.scala 12:21]
  wire  _T_981; // @[LZD.scala 49:16]
  wire  _T_982; // @[LZD.scala 49:27]
  wire  _T_983; // @[LZD.scala 49:25]
  wire [2:0] _T_984; // @[LZD.scala 49:47]
  wire [2:0] _T_985; // @[LZD.scala 49:59]
  wire [2:0] _T_986; // @[LZD.scala 49:35]
  wire [4:0] _T_988; // @[Cat.scala 29:58]
  wire [15:0] _T_989; // @[LZD.scala 44:32]
  wire [7:0] _T_990; // @[LZD.scala 43:32]
  wire [3:0] _T_991; // @[LZD.scala 43:32]
  wire [1:0] _T_992; // @[LZD.scala 43:32]
  wire  _T_993; // @[LZD.scala 39:14]
  wire  _T_994; // @[LZD.scala 39:21]
  wire  _T_995; // @[LZD.scala 39:30]
  wire  _T_996; // @[LZD.scala 39:27]
  wire  _T_997; // @[LZD.scala 39:25]
  wire [1:0] _T_998; // @[Cat.scala 29:58]
  wire [1:0] _T_999; // @[LZD.scala 44:32]
  wire  _T_1000; // @[LZD.scala 39:14]
  wire  _T_1001; // @[LZD.scala 39:21]
  wire  _T_1002; // @[LZD.scala 39:30]
  wire  _T_1003; // @[LZD.scala 39:27]
  wire  _T_1004; // @[LZD.scala 39:25]
  wire [1:0] _T_1005; // @[Cat.scala 29:58]
  wire  _T_1006; // @[Shift.scala 12:21]
  wire  _T_1007; // @[Shift.scala 12:21]
  wire  _T_1008; // @[LZD.scala 49:16]
  wire  _T_1009; // @[LZD.scala 49:27]
  wire  _T_1010; // @[LZD.scala 49:25]
  wire  _T_1011; // @[LZD.scala 49:47]
  wire  _T_1012; // @[LZD.scala 49:59]
  wire  _T_1013; // @[LZD.scala 49:35]
  wire [2:0] _T_1015; // @[Cat.scala 29:58]
  wire [3:0] _T_1016; // @[LZD.scala 44:32]
  wire [1:0] _T_1017; // @[LZD.scala 43:32]
  wire  _T_1018; // @[LZD.scala 39:14]
  wire  _T_1019; // @[LZD.scala 39:21]
  wire  _T_1020; // @[LZD.scala 39:30]
  wire  _T_1021; // @[LZD.scala 39:27]
  wire  _T_1022; // @[LZD.scala 39:25]
  wire [1:0] _T_1023; // @[Cat.scala 29:58]
  wire [1:0] _T_1024; // @[LZD.scala 44:32]
  wire  _T_1025; // @[LZD.scala 39:14]
  wire  _T_1026; // @[LZD.scala 39:21]
  wire  _T_1027; // @[LZD.scala 39:30]
  wire  _T_1028; // @[LZD.scala 39:27]
  wire  _T_1029; // @[LZD.scala 39:25]
  wire [1:0] _T_1030; // @[Cat.scala 29:58]
  wire  _T_1031; // @[Shift.scala 12:21]
  wire  _T_1032; // @[Shift.scala 12:21]
  wire  _T_1033; // @[LZD.scala 49:16]
  wire  _T_1034; // @[LZD.scala 49:27]
  wire  _T_1035; // @[LZD.scala 49:25]
  wire  _T_1036; // @[LZD.scala 49:47]
  wire  _T_1037; // @[LZD.scala 49:59]
  wire  _T_1038; // @[LZD.scala 49:35]
  wire [2:0] _T_1040; // @[Cat.scala 29:58]
  wire  _T_1041; // @[Shift.scala 12:21]
  wire  _T_1042; // @[Shift.scala 12:21]
  wire  _T_1043; // @[LZD.scala 49:16]
  wire  _T_1044; // @[LZD.scala 49:27]
  wire  _T_1045; // @[LZD.scala 49:25]
  wire [1:0] _T_1046; // @[LZD.scala 49:47]
  wire [1:0] _T_1047; // @[LZD.scala 49:59]
  wire [1:0] _T_1048; // @[LZD.scala 49:35]
  wire [3:0] _T_1050; // @[Cat.scala 29:58]
  wire [7:0] _T_1051; // @[LZD.scala 44:32]
  wire [3:0] _T_1052; // @[LZD.scala 43:32]
  wire [1:0] _T_1053; // @[LZD.scala 43:32]
  wire  _T_1054; // @[LZD.scala 39:14]
  wire  _T_1055; // @[LZD.scala 39:21]
  wire  _T_1056; // @[LZD.scala 39:30]
  wire  _T_1057; // @[LZD.scala 39:27]
  wire  _T_1058; // @[LZD.scala 39:25]
  wire [1:0] _T_1059; // @[Cat.scala 29:58]
  wire [1:0] _T_1060; // @[LZD.scala 44:32]
  wire  _T_1061; // @[LZD.scala 39:14]
  wire  _T_1062; // @[LZD.scala 39:21]
  wire  _T_1063; // @[LZD.scala 39:30]
  wire  _T_1064; // @[LZD.scala 39:27]
  wire  _T_1065; // @[LZD.scala 39:25]
  wire [1:0] _T_1066; // @[Cat.scala 29:58]
  wire  _T_1067; // @[Shift.scala 12:21]
  wire  _T_1068; // @[Shift.scala 12:21]
  wire  _T_1069; // @[LZD.scala 49:16]
  wire  _T_1070; // @[LZD.scala 49:27]
  wire  _T_1071; // @[LZD.scala 49:25]
  wire  _T_1072; // @[LZD.scala 49:47]
  wire  _T_1073; // @[LZD.scala 49:59]
  wire  _T_1074; // @[LZD.scala 49:35]
  wire [2:0] _T_1076; // @[Cat.scala 29:58]
  wire [3:0] _T_1077; // @[LZD.scala 44:32]
  wire [1:0] _T_1078; // @[LZD.scala 43:32]
  wire  _T_1079; // @[LZD.scala 39:14]
  wire  _T_1080; // @[LZD.scala 39:21]
  wire  _T_1081; // @[LZD.scala 39:30]
  wire  _T_1082; // @[LZD.scala 39:27]
  wire  _T_1083; // @[LZD.scala 39:25]
  wire [1:0] _T_1084; // @[Cat.scala 29:58]
  wire [1:0] _T_1085; // @[LZD.scala 44:32]
  wire  _T_1086; // @[LZD.scala 39:14]
  wire  _T_1087; // @[LZD.scala 39:21]
  wire  _T_1088; // @[LZD.scala 39:30]
  wire  _T_1089; // @[LZD.scala 39:27]
  wire  _T_1090; // @[LZD.scala 39:25]
  wire [1:0] _T_1091; // @[Cat.scala 29:58]
  wire  _T_1092; // @[Shift.scala 12:21]
  wire  _T_1093; // @[Shift.scala 12:21]
  wire  _T_1094; // @[LZD.scala 49:16]
  wire  _T_1095; // @[LZD.scala 49:27]
  wire  _T_1096; // @[LZD.scala 49:25]
  wire  _T_1097; // @[LZD.scala 49:47]
  wire  _T_1098; // @[LZD.scala 49:59]
  wire  _T_1099; // @[LZD.scala 49:35]
  wire [2:0] _T_1101; // @[Cat.scala 29:58]
  wire  _T_1102; // @[Shift.scala 12:21]
  wire  _T_1103; // @[Shift.scala 12:21]
  wire  _T_1104; // @[LZD.scala 49:16]
  wire  _T_1105; // @[LZD.scala 49:27]
  wire  _T_1106; // @[LZD.scala 49:25]
  wire [1:0] _T_1107; // @[LZD.scala 49:47]
  wire [1:0] _T_1108; // @[LZD.scala 49:59]
  wire [1:0] _T_1109; // @[LZD.scala 49:35]
  wire [3:0] _T_1111; // @[Cat.scala 29:58]
  wire  _T_1112; // @[Shift.scala 12:21]
  wire  _T_1113; // @[Shift.scala 12:21]
  wire  _T_1114; // @[LZD.scala 49:16]
  wire  _T_1115; // @[LZD.scala 49:27]
  wire  _T_1116; // @[LZD.scala 49:25]
  wire [2:0] _T_1117; // @[LZD.scala 49:47]
  wire [2:0] _T_1118; // @[LZD.scala 49:59]
  wire [2:0] _T_1119; // @[LZD.scala 49:35]
  wire [4:0] _T_1121; // @[Cat.scala 29:58]
  wire  _T_1122; // @[Shift.scala 12:21]
  wire  _T_1123; // @[Shift.scala 12:21]
  wire  _T_1124; // @[LZD.scala 49:16]
  wire  _T_1125; // @[LZD.scala 49:27]
  wire  _T_1126; // @[LZD.scala 49:25]
  wire [3:0] _T_1127; // @[LZD.scala 49:47]
  wire [3:0] _T_1128; // @[LZD.scala 49:59]
  wire [3:0] _T_1129; // @[LZD.scala 49:35]
  wire [5:0] _T_1131; // @[Cat.scala 29:58]
  wire  _T_1132; // @[Shift.scala 12:21]
  wire  _T_1133; // @[Shift.scala 12:21]
  wire  _T_1134; // @[LZD.scala 49:16]
  wire  _T_1135; // @[LZD.scala 49:27]
  wire  _T_1136; // @[LZD.scala 49:25]
  wire [4:0] _T_1137; // @[LZD.scala 49:47]
  wire [4:0] _T_1138; // @[LZD.scala 49:59]
  wire [4:0] _T_1139; // @[LZD.scala 49:35]
  wire [6:0] _T_1141; // @[Cat.scala 29:58]
  wire  _T_1142; // @[Shift.scala 12:21]
  wire  _T_1143; // @[Shift.scala 12:21]
  wire  _T_1144; // @[LZD.scala 49:16]
  wire  _T_1145; // @[LZD.scala 49:27]
  wire  _T_1146; // @[LZD.scala 49:25]
  wire [5:0] _T_1147; // @[LZD.scala 49:47]
  wire [5:0] _T_1148; // @[LZD.scala 49:59]
  wire [5:0] _T_1149; // @[LZD.scala 49:35]
  wire [7:0] _T_1151; // @[Cat.scala 29:58]
  wire [127:0] _T_1152; // @[LZD.scala 44:32]
  wire [63:0] _T_1153; // @[LZD.scala 43:32]
  wire [31:0] _T_1154; // @[LZD.scala 43:32]
  wire [15:0] _T_1155; // @[LZD.scala 43:32]
  wire [7:0] _T_1156; // @[LZD.scala 43:32]
  wire [3:0] _T_1157; // @[LZD.scala 43:32]
  wire [1:0] _T_1158; // @[LZD.scala 43:32]
  wire  _T_1159; // @[LZD.scala 39:14]
  wire  _T_1160; // @[LZD.scala 39:21]
  wire  _T_1161; // @[LZD.scala 39:30]
  wire  _T_1162; // @[LZD.scala 39:27]
  wire  _T_1163; // @[LZD.scala 39:25]
  wire [1:0] _T_1164; // @[Cat.scala 29:58]
  wire [1:0] _T_1165; // @[LZD.scala 44:32]
  wire  _T_1166; // @[LZD.scala 39:14]
  wire  _T_1167; // @[LZD.scala 39:21]
  wire  _T_1168; // @[LZD.scala 39:30]
  wire  _T_1169; // @[LZD.scala 39:27]
  wire  _T_1170; // @[LZD.scala 39:25]
  wire [1:0] _T_1171; // @[Cat.scala 29:58]
  wire  _T_1172; // @[Shift.scala 12:21]
  wire  _T_1173; // @[Shift.scala 12:21]
  wire  _T_1174; // @[LZD.scala 49:16]
  wire  _T_1175; // @[LZD.scala 49:27]
  wire  _T_1176; // @[LZD.scala 49:25]
  wire  _T_1177; // @[LZD.scala 49:47]
  wire  _T_1178; // @[LZD.scala 49:59]
  wire  _T_1179; // @[LZD.scala 49:35]
  wire [2:0] _T_1181; // @[Cat.scala 29:58]
  wire [3:0] _T_1182; // @[LZD.scala 44:32]
  wire [1:0] _T_1183; // @[LZD.scala 43:32]
  wire  _T_1184; // @[LZD.scala 39:14]
  wire  _T_1185; // @[LZD.scala 39:21]
  wire  _T_1186; // @[LZD.scala 39:30]
  wire  _T_1187; // @[LZD.scala 39:27]
  wire  _T_1188; // @[LZD.scala 39:25]
  wire [1:0] _T_1189; // @[Cat.scala 29:58]
  wire [1:0] _T_1190; // @[LZD.scala 44:32]
  wire  _T_1191; // @[LZD.scala 39:14]
  wire  _T_1192; // @[LZD.scala 39:21]
  wire  _T_1193; // @[LZD.scala 39:30]
  wire  _T_1194; // @[LZD.scala 39:27]
  wire  _T_1195; // @[LZD.scala 39:25]
  wire [1:0] _T_1196; // @[Cat.scala 29:58]
  wire  _T_1197; // @[Shift.scala 12:21]
  wire  _T_1198; // @[Shift.scala 12:21]
  wire  _T_1199; // @[LZD.scala 49:16]
  wire  _T_1200; // @[LZD.scala 49:27]
  wire  _T_1201; // @[LZD.scala 49:25]
  wire  _T_1202; // @[LZD.scala 49:47]
  wire  _T_1203; // @[LZD.scala 49:59]
  wire  _T_1204; // @[LZD.scala 49:35]
  wire [2:0] _T_1206; // @[Cat.scala 29:58]
  wire  _T_1207; // @[Shift.scala 12:21]
  wire  _T_1208; // @[Shift.scala 12:21]
  wire  _T_1209; // @[LZD.scala 49:16]
  wire  _T_1210; // @[LZD.scala 49:27]
  wire  _T_1211; // @[LZD.scala 49:25]
  wire [1:0] _T_1212; // @[LZD.scala 49:47]
  wire [1:0] _T_1213; // @[LZD.scala 49:59]
  wire [1:0] _T_1214; // @[LZD.scala 49:35]
  wire [3:0] _T_1216; // @[Cat.scala 29:58]
  wire [7:0] _T_1217; // @[LZD.scala 44:32]
  wire [3:0] _T_1218; // @[LZD.scala 43:32]
  wire [1:0] _T_1219; // @[LZD.scala 43:32]
  wire  _T_1220; // @[LZD.scala 39:14]
  wire  _T_1221; // @[LZD.scala 39:21]
  wire  _T_1222; // @[LZD.scala 39:30]
  wire  _T_1223; // @[LZD.scala 39:27]
  wire  _T_1224; // @[LZD.scala 39:25]
  wire [1:0] _T_1225; // @[Cat.scala 29:58]
  wire [1:0] _T_1226; // @[LZD.scala 44:32]
  wire  _T_1227; // @[LZD.scala 39:14]
  wire  _T_1228; // @[LZD.scala 39:21]
  wire  _T_1229; // @[LZD.scala 39:30]
  wire  _T_1230; // @[LZD.scala 39:27]
  wire  _T_1231; // @[LZD.scala 39:25]
  wire [1:0] _T_1232; // @[Cat.scala 29:58]
  wire  _T_1233; // @[Shift.scala 12:21]
  wire  _T_1234; // @[Shift.scala 12:21]
  wire  _T_1235; // @[LZD.scala 49:16]
  wire  _T_1236; // @[LZD.scala 49:27]
  wire  _T_1237; // @[LZD.scala 49:25]
  wire  _T_1238; // @[LZD.scala 49:47]
  wire  _T_1239; // @[LZD.scala 49:59]
  wire  _T_1240; // @[LZD.scala 49:35]
  wire [2:0] _T_1242; // @[Cat.scala 29:58]
  wire [3:0] _T_1243; // @[LZD.scala 44:32]
  wire [1:0] _T_1244; // @[LZD.scala 43:32]
  wire  _T_1245; // @[LZD.scala 39:14]
  wire  _T_1246; // @[LZD.scala 39:21]
  wire  _T_1247; // @[LZD.scala 39:30]
  wire  _T_1248; // @[LZD.scala 39:27]
  wire  _T_1249; // @[LZD.scala 39:25]
  wire [1:0] _T_1250; // @[Cat.scala 29:58]
  wire [1:0] _T_1251; // @[LZD.scala 44:32]
  wire  _T_1252; // @[LZD.scala 39:14]
  wire  _T_1253; // @[LZD.scala 39:21]
  wire  _T_1254; // @[LZD.scala 39:30]
  wire  _T_1255; // @[LZD.scala 39:27]
  wire  _T_1256; // @[LZD.scala 39:25]
  wire [1:0] _T_1257; // @[Cat.scala 29:58]
  wire  _T_1258; // @[Shift.scala 12:21]
  wire  _T_1259; // @[Shift.scala 12:21]
  wire  _T_1260; // @[LZD.scala 49:16]
  wire  _T_1261; // @[LZD.scala 49:27]
  wire  _T_1262; // @[LZD.scala 49:25]
  wire  _T_1263; // @[LZD.scala 49:47]
  wire  _T_1264; // @[LZD.scala 49:59]
  wire  _T_1265; // @[LZD.scala 49:35]
  wire [2:0] _T_1267; // @[Cat.scala 29:58]
  wire  _T_1268; // @[Shift.scala 12:21]
  wire  _T_1269; // @[Shift.scala 12:21]
  wire  _T_1270; // @[LZD.scala 49:16]
  wire  _T_1271; // @[LZD.scala 49:27]
  wire  _T_1272; // @[LZD.scala 49:25]
  wire [1:0] _T_1273; // @[LZD.scala 49:47]
  wire [1:0] _T_1274; // @[LZD.scala 49:59]
  wire [1:0] _T_1275; // @[LZD.scala 49:35]
  wire [3:0] _T_1277; // @[Cat.scala 29:58]
  wire  _T_1278; // @[Shift.scala 12:21]
  wire  _T_1279; // @[Shift.scala 12:21]
  wire  _T_1280; // @[LZD.scala 49:16]
  wire  _T_1281; // @[LZD.scala 49:27]
  wire  _T_1282; // @[LZD.scala 49:25]
  wire [2:0] _T_1283; // @[LZD.scala 49:47]
  wire [2:0] _T_1284; // @[LZD.scala 49:59]
  wire [2:0] _T_1285; // @[LZD.scala 49:35]
  wire [4:0] _T_1287; // @[Cat.scala 29:58]
  wire [15:0] _T_1288; // @[LZD.scala 44:32]
  wire [7:0] _T_1289; // @[LZD.scala 43:32]
  wire [3:0] _T_1290; // @[LZD.scala 43:32]
  wire [1:0] _T_1291; // @[LZD.scala 43:32]
  wire  _T_1292; // @[LZD.scala 39:14]
  wire  _T_1293; // @[LZD.scala 39:21]
  wire  _T_1294; // @[LZD.scala 39:30]
  wire  _T_1295; // @[LZD.scala 39:27]
  wire  _T_1296; // @[LZD.scala 39:25]
  wire [1:0] _T_1297; // @[Cat.scala 29:58]
  wire [1:0] _T_1298; // @[LZD.scala 44:32]
  wire  _T_1299; // @[LZD.scala 39:14]
  wire  _T_1300; // @[LZD.scala 39:21]
  wire  _T_1301; // @[LZD.scala 39:30]
  wire  _T_1302; // @[LZD.scala 39:27]
  wire  _T_1303; // @[LZD.scala 39:25]
  wire [1:0] _T_1304; // @[Cat.scala 29:58]
  wire  _T_1305; // @[Shift.scala 12:21]
  wire  _T_1306; // @[Shift.scala 12:21]
  wire  _T_1307; // @[LZD.scala 49:16]
  wire  _T_1308; // @[LZD.scala 49:27]
  wire  _T_1309; // @[LZD.scala 49:25]
  wire  _T_1310; // @[LZD.scala 49:47]
  wire  _T_1311; // @[LZD.scala 49:59]
  wire  _T_1312; // @[LZD.scala 49:35]
  wire [2:0] _T_1314; // @[Cat.scala 29:58]
  wire [3:0] _T_1315; // @[LZD.scala 44:32]
  wire [1:0] _T_1316; // @[LZD.scala 43:32]
  wire  _T_1317; // @[LZD.scala 39:14]
  wire  _T_1318; // @[LZD.scala 39:21]
  wire  _T_1319; // @[LZD.scala 39:30]
  wire  _T_1320; // @[LZD.scala 39:27]
  wire  _T_1321; // @[LZD.scala 39:25]
  wire [1:0] _T_1322; // @[Cat.scala 29:58]
  wire [1:0] _T_1323; // @[LZD.scala 44:32]
  wire  _T_1324; // @[LZD.scala 39:14]
  wire  _T_1325; // @[LZD.scala 39:21]
  wire  _T_1326; // @[LZD.scala 39:30]
  wire  _T_1327; // @[LZD.scala 39:27]
  wire  _T_1328; // @[LZD.scala 39:25]
  wire [1:0] _T_1329; // @[Cat.scala 29:58]
  wire  _T_1330; // @[Shift.scala 12:21]
  wire  _T_1331; // @[Shift.scala 12:21]
  wire  _T_1332; // @[LZD.scala 49:16]
  wire  _T_1333; // @[LZD.scala 49:27]
  wire  _T_1334; // @[LZD.scala 49:25]
  wire  _T_1335; // @[LZD.scala 49:47]
  wire  _T_1336; // @[LZD.scala 49:59]
  wire  _T_1337; // @[LZD.scala 49:35]
  wire [2:0] _T_1339; // @[Cat.scala 29:58]
  wire  _T_1340; // @[Shift.scala 12:21]
  wire  _T_1341; // @[Shift.scala 12:21]
  wire  _T_1342; // @[LZD.scala 49:16]
  wire  _T_1343; // @[LZD.scala 49:27]
  wire  _T_1344; // @[LZD.scala 49:25]
  wire [1:0] _T_1345; // @[LZD.scala 49:47]
  wire [1:0] _T_1346; // @[LZD.scala 49:59]
  wire [1:0] _T_1347; // @[LZD.scala 49:35]
  wire [3:0] _T_1349; // @[Cat.scala 29:58]
  wire [7:0] _T_1350; // @[LZD.scala 44:32]
  wire [3:0] _T_1351; // @[LZD.scala 43:32]
  wire [1:0] _T_1352; // @[LZD.scala 43:32]
  wire  _T_1353; // @[LZD.scala 39:14]
  wire  _T_1354; // @[LZD.scala 39:21]
  wire  _T_1355; // @[LZD.scala 39:30]
  wire  _T_1356; // @[LZD.scala 39:27]
  wire  _T_1357; // @[LZD.scala 39:25]
  wire [1:0] _T_1358; // @[Cat.scala 29:58]
  wire [1:0] _T_1359; // @[LZD.scala 44:32]
  wire  _T_1360; // @[LZD.scala 39:14]
  wire  _T_1361; // @[LZD.scala 39:21]
  wire  _T_1362; // @[LZD.scala 39:30]
  wire  _T_1363; // @[LZD.scala 39:27]
  wire  _T_1364; // @[LZD.scala 39:25]
  wire [1:0] _T_1365; // @[Cat.scala 29:58]
  wire  _T_1366; // @[Shift.scala 12:21]
  wire  _T_1367; // @[Shift.scala 12:21]
  wire  _T_1368; // @[LZD.scala 49:16]
  wire  _T_1369; // @[LZD.scala 49:27]
  wire  _T_1370; // @[LZD.scala 49:25]
  wire  _T_1371; // @[LZD.scala 49:47]
  wire  _T_1372; // @[LZD.scala 49:59]
  wire  _T_1373; // @[LZD.scala 49:35]
  wire [2:0] _T_1375; // @[Cat.scala 29:58]
  wire [3:0] _T_1376; // @[LZD.scala 44:32]
  wire [1:0] _T_1377; // @[LZD.scala 43:32]
  wire  _T_1378; // @[LZD.scala 39:14]
  wire  _T_1379; // @[LZD.scala 39:21]
  wire  _T_1380; // @[LZD.scala 39:30]
  wire  _T_1381; // @[LZD.scala 39:27]
  wire  _T_1382; // @[LZD.scala 39:25]
  wire [1:0] _T_1383; // @[Cat.scala 29:58]
  wire [1:0] _T_1384; // @[LZD.scala 44:32]
  wire  _T_1385; // @[LZD.scala 39:14]
  wire  _T_1386; // @[LZD.scala 39:21]
  wire  _T_1387; // @[LZD.scala 39:30]
  wire  _T_1388; // @[LZD.scala 39:27]
  wire  _T_1389; // @[LZD.scala 39:25]
  wire [1:0] _T_1390; // @[Cat.scala 29:58]
  wire  _T_1391; // @[Shift.scala 12:21]
  wire  _T_1392; // @[Shift.scala 12:21]
  wire  _T_1393; // @[LZD.scala 49:16]
  wire  _T_1394; // @[LZD.scala 49:27]
  wire  _T_1395; // @[LZD.scala 49:25]
  wire  _T_1396; // @[LZD.scala 49:47]
  wire  _T_1397; // @[LZD.scala 49:59]
  wire  _T_1398; // @[LZD.scala 49:35]
  wire [2:0] _T_1400; // @[Cat.scala 29:58]
  wire  _T_1401; // @[Shift.scala 12:21]
  wire  _T_1402; // @[Shift.scala 12:21]
  wire  _T_1403; // @[LZD.scala 49:16]
  wire  _T_1404; // @[LZD.scala 49:27]
  wire  _T_1405; // @[LZD.scala 49:25]
  wire [1:0] _T_1406; // @[LZD.scala 49:47]
  wire [1:0] _T_1407; // @[LZD.scala 49:59]
  wire [1:0] _T_1408; // @[LZD.scala 49:35]
  wire [3:0] _T_1410; // @[Cat.scala 29:58]
  wire  _T_1411; // @[Shift.scala 12:21]
  wire  _T_1412; // @[Shift.scala 12:21]
  wire  _T_1413; // @[LZD.scala 49:16]
  wire  _T_1414; // @[LZD.scala 49:27]
  wire  _T_1415; // @[LZD.scala 49:25]
  wire [2:0] _T_1416; // @[LZD.scala 49:47]
  wire [2:0] _T_1417; // @[LZD.scala 49:59]
  wire [2:0] _T_1418; // @[LZD.scala 49:35]
  wire [4:0] _T_1420; // @[Cat.scala 29:58]
  wire  _T_1421; // @[Shift.scala 12:21]
  wire  _T_1422; // @[Shift.scala 12:21]
  wire  _T_1423; // @[LZD.scala 49:16]
  wire  _T_1424; // @[LZD.scala 49:27]
  wire  _T_1425; // @[LZD.scala 49:25]
  wire [3:0] _T_1426; // @[LZD.scala 49:47]
  wire [3:0] _T_1427; // @[LZD.scala 49:59]
  wire [3:0] _T_1428; // @[LZD.scala 49:35]
  wire [5:0] _T_1430; // @[Cat.scala 29:58]
  wire [31:0] _T_1431; // @[LZD.scala 44:32]
  wire [15:0] _T_1432; // @[LZD.scala 43:32]
  wire [7:0] _T_1433; // @[LZD.scala 43:32]
  wire [3:0] _T_1434; // @[LZD.scala 43:32]
  wire [1:0] _T_1435; // @[LZD.scala 43:32]
  wire  _T_1436; // @[LZD.scala 39:14]
  wire  _T_1437; // @[LZD.scala 39:21]
  wire  _T_1438; // @[LZD.scala 39:30]
  wire  _T_1439; // @[LZD.scala 39:27]
  wire  _T_1440; // @[LZD.scala 39:25]
  wire [1:0] _T_1441; // @[Cat.scala 29:58]
  wire [1:0] _T_1442; // @[LZD.scala 44:32]
  wire  _T_1443; // @[LZD.scala 39:14]
  wire  _T_1444; // @[LZD.scala 39:21]
  wire  _T_1445; // @[LZD.scala 39:30]
  wire  _T_1446; // @[LZD.scala 39:27]
  wire  _T_1447; // @[LZD.scala 39:25]
  wire [1:0] _T_1448; // @[Cat.scala 29:58]
  wire  _T_1449; // @[Shift.scala 12:21]
  wire  _T_1450; // @[Shift.scala 12:21]
  wire  _T_1451; // @[LZD.scala 49:16]
  wire  _T_1452; // @[LZD.scala 49:27]
  wire  _T_1453; // @[LZD.scala 49:25]
  wire  _T_1454; // @[LZD.scala 49:47]
  wire  _T_1455; // @[LZD.scala 49:59]
  wire  _T_1456; // @[LZD.scala 49:35]
  wire [2:0] _T_1458; // @[Cat.scala 29:58]
  wire [3:0] _T_1459; // @[LZD.scala 44:32]
  wire [1:0] _T_1460; // @[LZD.scala 43:32]
  wire  _T_1461; // @[LZD.scala 39:14]
  wire  _T_1462; // @[LZD.scala 39:21]
  wire  _T_1463; // @[LZD.scala 39:30]
  wire  _T_1464; // @[LZD.scala 39:27]
  wire  _T_1465; // @[LZD.scala 39:25]
  wire [1:0] _T_1466; // @[Cat.scala 29:58]
  wire [1:0] _T_1467; // @[LZD.scala 44:32]
  wire  _T_1468; // @[LZD.scala 39:14]
  wire  _T_1469; // @[LZD.scala 39:21]
  wire  _T_1470; // @[LZD.scala 39:30]
  wire  _T_1471; // @[LZD.scala 39:27]
  wire  _T_1472; // @[LZD.scala 39:25]
  wire [1:0] _T_1473; // @[Cat.scala 29:58]
  wire  _T_1474; // @[Shift.scala 12:21]
  wire  _T_1475; // @[Shift.scala 12:21]
  wire  _T_1476; // @[LZD.scala 49:16]
  wire  _T_1477; // @[LZD.scala 49:27]
  wire  _T_1478; // @[LZD.scala 49:25]
  wire  _T_1479; // @[LZD.scala 49:47]
  wire  _T_1480; // @[LZD.scala 49:59]
  wire  _T_1481; // @[LZD.scala 49:35]
  wire [2:0] _T_1483; // @[Cat.scala 29:58]
  wire  _T_1484; // @[Shift.scala 12:21]
  wire  _T_1485; // @[Shift.scala 12:21]
  wire  _T_1486; // @[LZD.scala 49:16]
  wire  _T_1487; // @[LZD.scala 49:27]
  wire  _T_1488; // @[LZD.scala 49:25]
  wire [1:0] _T_1489; // @[LZD.scala 49:47]
  wire [1:0] _T_1490; // @[LZD.scala 49:59]
  wire [1:0] _T_1491; // @[LZD.scala 49:35]
  wire [3:0] _T_1493; // @[Cat.scala 29:58]
  wire [7:0] _T_1494; // @[LZD.scala 44:32]
  wire [3:0] _T_1495; // @[LZD.scala 43:32]
  wire [1:0] _T_1496; // @[LZD.scala 43:32]
  wire  _T_1497; // @[LZD.scala 39:14]
  wire  _T_1498; // @[LZD.scala 39:21]
  wire  _T_1499; // @[LZD.scala 39:30]
  wire  _T_1500; // @[LZD.scala 39:27]
  wire  _T_1501; // @[LZD.scala 39:25]
  wire [1:0] _T_1502; // @[Cat.scala 29:58]
  wire [1:0] _T_1503; // @[LZD.scala 44:32]
  wire  _T_1504; // @[LZD.scala 39:14]
  wire  _T_1505; // @[LZD.scala 39:21]
  wire  _T_1506; // @[LZD.scala 39:30]
  wire  _T_1507; // @[LZD.scala 39:27]
  wire  _T_1508; // @[LZD.scala 39:25]
  wire [1:0] _T_1509; // @[Cat.scala 29:58]
  wire  _T_1510; // @[Shift.scala 12:21]
  wire  _T_1511; // @[Shift.scala 12:21]
  wire  _T_1512; // @[LZD.scala 49:16]
  wire  _T_1513; // @[LZD.scala 49:27]
  wire  _T_1514; // @[LZD.scala 49:25]
  wire  _T_1515; // @[LZD.scala 49:47]
  wire  _T_1516; // @[LZD.scala 49:59]
  wire  _T_1517; // @[LZD.scala 49:35]
  wire [2:0] _T_1519; // @[Cat.scala 29:58]
  wire [3:0] _T_1520; // @[LZD.scala 44:32]
  wire [1:0] _T_1521; // @[LZD.scala 43:32]
  wire  _T_1522; // @[LZD.scala 39:14]
  wire  _T_1523; // @[LZD.scala 39:21]
  wire  _T_1524; // @[LZD.scala 39:30]
  wire  _T_1525; // @[LZD.scala 39:27]
  wire  _T_1526; // @[LZD.scala 39:25]
  wire [1:0] _T_1527; // @[Cat.scala 29:58]
  wire [1:0] _T_1528; // @[LZD.scala 44:32]
  wire  _T_1529; // @[LZD.scala 39:14]
  wire  _T_1530; // @[LZD.scala 39:21]
  wire  _T_1531; // @[LZD.scala 39:30]
  wire  _T_1532; // @[LZD.scala 39:27]
  wire  _T_1533; // @[LZD.scala 39:25]
  wire [1:0] _T_1534; // @[Cat.scala 29:58]
  wire  _T_1535; // @[Shift.scala 12:21]
  wire  _T_1536; // @[Shift.scala 12:21]
  wire  _T_1537; // @[LZD.scala 49:16]
  wire  _T_1538; // @[LZD.scala 49:27]
  wire  _T_1539; // @[LZD.scala 49:25]
  wire  _T_1540; // @[LZD.scala 49:47]
  wire  _T_1541; // @[LZD.scala 49:59]
  wire  _T_1542; // @[LZD.scala 49:35]
  wire [2:0] _T_1544; // @[Cat.scala 29:58]
  wire  _T_1545; // @[Shift.scala 12:21]
  wire  _T_1546; // @[Shift.scala 12:21]
  wire  _T_1547; // @[LZD.scala 49:16]
  wire  _T_1548; // @[LZD.scala 49:27]
  wire  _T_1549; // @[LZD.scala 49:25]
  wire [1:0] _T_1550; // @[LZD.scala 49:47]
  wire [1:0] _T_1551; // @[LZD.scala 49:59]
  wire [1:0] _T_1552; // @[LZD.scala 49:35]
  wire [3:0] _T_1554; // @[Cat.scala 29:58]
  wire  _T_1555; // @[Shift.scala 12:21]
  wire  _T_1556; // @[Shift.scala 12:21]
  wire  _T_1557; // @[LZD.scala 49:16]
  wire  _T_1558; // @[LZD.scala 49:27]
  wire  _T_1559; // @[LZD.scala 49:25]
  wire [2:0] _T_1560; // @[LZD.scala 49:47]
  wire [2:0] _T_1561; // @[LZD.scala 49:59]
  wire [2:0] _T_1562; // @[LZD.scala 49:35]
  wire [4:0] _T_1564; // @[Cat.scala 29:58]
  wire [15:0] _T_1565; // @[LZD.scala 44:32]
  wire [7:0] _T_1566; // @[LZD.scala 43:32]
  wire [3:0] _T_1567; // @[LZD.scala 43:32]
  wire [1:0] _T_1568; // @[LZD.scala 43:32]
  wire  _T_1569; // @[LZD.scala 39:14]
  wire  _T_1570; // @[LZD.scala 39:21]
  wire  _T_1571; // @[LZD.scala 39:30]
  wire  _T_1572; // @[LZD.scala 39:27]
  wire  _T_1573; // @[LZD.scala 39:25]
  wire [1:0] _T_1574; // @[Cat.scala 29:58]
  wire [1:0] _T_1575; // @[LZD.scala 44:32]
  wire  _T_1576; // @[LZD.scala 39:14]
  wire  _T_1577; // @[LZD.scala 39:21]
  wire  _T_1578; // @[LZD.scala 39:30]
  wire  _T_1579; // @[LZD.scala 39:27]
  wire  _T_1580; // @[LZD.scala 39:25]
  wire [1:0] _T_1581; // @[Cat.scala 29:58]
  wire  _T_1582; // @[Shift.scala 12:21]
  wire  _T_1583; // @[Shift.scala 12:21]
  wire  _T_1584; // @[LZD.scala 49:16]
  wire  _T_1585; // @[LZD.scala 49:27]
  wire  _T_1586; // @[LZD.scala 49:25]
  wire  _T_1587; // @[LZD.scala 49:47]
  wire  _T_1588; // @[LZD.scala 49:59]
  wire  _T_1589; // @[LZD.scala 49:35]
  wire [2:0] _T_1591; // @[Cat.scala 29:58]
  wire [3:0] _T_1592; // @[LZD.scala 44:32]
  wire [1:0] _T_1593; // @[LZD.scala 43:32]
  wire  _T_1594; // @[LZD.scala 39:14]
  wire  _T_1595; // @[LZD.scala 39:21]
  wire  _T_1596; // @[LZD.scala 39:30]
  wire  _T_1597; // @[LZD.scala 39:27]
  wire  _T_1598; // @[LZD.scala 39:25]
  wire [1:0] _T_1599; // @[Cat.scala 29:58]
  wire [1:0] _T_1600; // @[LZD.scala 44:32]
  wire  _T_1601; // @[LZD.scala 39:14]
  wire  _T_1602; // @[LZD.scala 39:21]
  wire  _T_1603; // @[LZD.scala 39:30]
  wire  _T_1604; // @[LZD.scala 39:27]
  wire  _T_1605; // @[LZD.scala 39:25]
  wire [1:0] _T_1606; // @[Cat.scala 29:58]
  wire  _T_1607; // @[Shift.scala 12:21]
  wire  _T_1608; // @[Shift.scala 12:21]
  wire  _T_1609; // @[LZD.scala 49:16]
  wire  _T_1610; // @[LZD.scala 49:27]
  wire  _T_1611; // @[LZD.scala 49:25]
  wire  _T_1612; // @[LZD.scala 49:47]
  wire  _T_1613; // @[LZD.scala 49:59]
  wire  _T_1614; // @[LZD.scala 49:35]
  wire [2:0] _T_1616; // @[Cat.scala 29:58]
  wire  _T_1617; // @[Shift.scala 12:21]
  wire  _T_1618; // @[Shift.scala 12:21]
  wire  _T_1619; // @[LZD.scala 49:16]
  wire  _T_1620; // @[LZD.scala 49:27]
  wire  _T_1621; // @[LZD.scala 49:25]
  wire [1:0] _T_1622; // @[LZD.scala 49:47]
  wire [1:0] _T_1623; // @[LZD.scala 49:59]
  wire [1:0] _T_1624; // @[LZD.scala 49:35]
  wire [3:0] _T_1626; // @[Cat.scala 29:58]
  wire [7:0] _T_1627; // @[LZD.scala 44:32]
  wire [3:0] _T_1628; // @[LZD.scala 43:32]
  wire [1:0] _T_1629; // @[LZD.scala 43:32]
  wire  _T_1630; // @[LZD.scala 39:14]
  wire  _T_1631; // @[LZD.scala 39:21]
  wire  _T_1632; // @[LZD.scala 39:30]
  wire  _T_1633; // @[LZD.scala 39:27]
  wire  _T_1634; // @[LZD.scala 39:25]
  wire [1:0] _T_1635; // @[Cat.scala 29:58]
  wire [1:0] _T_1636; // @[LZD.scala 44:32]
  wire  _T_1637; // @[LZD.scala 39:14]
  wire  _T_1638; // @[LZD.scala 39:21]
  wire  _T_1639; // @[LZD.scala 39:30]
  wire  _T_1640; // @[LZD.scala 39:27]
  wire  _T_1641; // @[LZD.scala 39:25]
  wire [1:0] _T_1642; // @[Cat.scala 29:58]
  wire  _T_1643; // @[Shift.scala 12:21]
  wire  _T_1644; // @[Shift.scala 12:21]
  wire  _T_1645; // @[LZD.scala 49:16]
  wire  _T_1646; // @[LZD.scala 49:27]
  wire  _T_1647; // @[LZD.scala 49:25]
  wire  _T_1648; // @[LZD.scala 49:47]
  wire  _T_1649; // @[LZD.scala 49:59]
  wire  _T_1650; // @[LZD.scala 49:35]
  wire [2:0] _T_1652; // @[Cat.scala 29:58]
  wire [3:0] _T_1653; // @[LZD.scala 44:32]
  wire [1:0] _T_1654; // @[LZD.scala 43:32]
  wire  _T_1655; // @[LZD.scala 39:14]
  wire  _T_1656; // @[LZD.scala 39:21]
  wire  _T_1657; // @[LZD.scala 39:30]
  wire  _T_1658; // @[LZD.scala 39:27]
  wire  _T_1659; // @[LZD.scala 39:25]
  wire [1:0] _T_1660; // @[Cat.scala 29:58]
  wire [1:0] _T_1661; // @[LZD.scala 44:32]
  wire  _T_1662; // @[LZD.scala 39:14]
  wire  _T_1663; // @[LZD.scala 39:21]
  wire  _T_1664; // @[LZD.scala 39:30]
  wire  _T_1665; // @[LZD.scala 39:27]
  wire  _T_1666; // @[LZD.scala 39:25]
  wire [1:0] _T_1667; // @[Cat.scala 29:58]
  wire  _T_1668; // @[Shift.scala 12:21]
  wire  _T_1669; // @[Shift.scala 12:21]
  wire  _T_1670; // @[LZD.scala 49:16]
  wire  _T_1671; // @[LZD.scala 49:27]
  wire  _T_1672; // @[LZD.scala 49:25]
  wire  _T_1673; // @[LZD.scala 49:47]
  wire  _T_1674; // @[LZD.scala 49:59]
  wire  _T_1675; // @[LZD.scala 49:35]
  wire [2:0] _T_1677; // @[Cat.scala 29:58]
  wire  _T_1678; // @[Shift.scala 12:21]
  wire  _T_1679; // @[Shift.scala 12:21]
  wire  _T_1680; // @[LZD.scala 49:16]
  wire  _T_1681; // @[LZD.scala 49:27]
  wire  _T_1682; // @[LZD.scala 49:25]
  wire [1:0] _T_1683; // @[LZD.scala 49:47]
  wire [1:0] _T_1684; // @[LZD.scala 49:59]
  wire [1:0] _T_1685; // @[LZD.scala 49:35]
  wire [3:0] _T_1687; // @[Cat.scala 29:58]
  wire  _T_1688; // @[Shift.scala 12:21]
  wire  _T_1689; // @[Shift.scala 12:21]
  wire  _T_1690; // @[LZD.scala 49:16]
  wire  _T_1691; // @[LZD.scala 49:27]
  wire  _T_1692; // @[LZD.scala 49:25]
  wire [2:0] _T_1693; // @[LZD.scala 49:47]
  wire [2:0] _T_1694; // @[LZD.scala 49:59]
  wire [2:0] _T_1695; // @[LZD.scala 49:35]
  wire [4:0] _T_1697; // @[Cat.scala 29:58]
  wire  _T_1698; // @[Shift.scala 12:21]
  wire  _T_1699; // @[Shift.scala 12:21]
  wire  _T_1700; // @[LZD.scala 49:16]
  wire  _T_1701; // @[LZD.scala 49:27]
  wire  _T_1702; // @[LZD.scala 49:25]
  wire [3:0] _T_1703; // @[LZD.scala 49:47]
  wire [3:0] _T_1704; // @[LZD.scala 49:59]
  wire [3:0] _T_1705; // @[LZD.scala 49:35]
  wire [5:0] _T_1707; // @[Cat.scala 29:58]
  wire  _T_1708; // @[Shift.scala 12:21]
  wire  _T_1709; // @[Shift.scala 12:21]
  wire  _T_1710; // @[LZD.scala 49:16]
  wire  _T_1711; // @[LZD.scala 49:27]
  wire  _T_1712; // @[LZD.scala 49:25]
  wire [4:0] _T_1713; // @[LZD.scala 49:47]
  wire [4:0] _T_1714; // @[LZD.scala 49:59]
  wire [4:0] _T_1715; // @[LZD.scala 49:35]
  wire [6:0] _T_1717; // @[Cat.scala 29:58]
  wire [63:0] _T_1718; // @[LZD.scala 44:32]
  wire [31:0] _T_1719; // @[LZD.scala 43:32]
  wire [15:0] _T_1720; // @[LZD.scala 43:32]
  wire [7:0] _T_1721; // @[LZD.scala 43:32]
  wire [3:0] _T_1722; // @[LZD.scala 43:32]
  wire [1:0] _T_1723; // @[LZD.scala 43:32]
  wire  _T_1724; // @[LZD.scala 39:14]
  wire  _T_1725; // @[LZD.scala 39:21]
  wire  _T_1726; // @[LZD.scala 39:30]
  wire  _T_1727; // @[LZD.scala 39:27]
  wire  _T_1728; // @[LZD.scala 39:25]
  wire [1:0] _T_1729; // @[Cat.scala 29:58]
  wire [1:0] _T_1730; // @[LZD.scala 44:32]
  wire  _T_1731; // @[LZD.scala 39:14]
  wire  _T_1732; // @[LZD.scala 39:21]
  wire  _T_1733; // @[LZD.scala 39:30]
  wire  _T_1734; // @[LZD.scala 39:27]
  wire  _T_1735; // @[LZD.scala 39:25]
  wire [1:0] _T_1736; // @[Cat.scala 29:58]
  wire  _T_1737; // @[Shift.scala 12:21]
  wire  _T_1738; // @[Shift.scala 12:21]
  wire  _T_1739; // @[LZD.scala 49:16]
  wire  _T_1740; // @[LZD.scala 49:27]
  wire  _T_1741; // @[LZD.scala 49:25]
  wire  _T_1742; // @[LZD.scala 49:47]
  wire  _T_1743; // @[LZD.scala 49:59]
  wire  _T_1744; // @[LZD.scala 49:35]
  wire [2:0] _T_1746; // @[Cat.scala 29:58]
  wire [3:0] _T_1747; // @[LZD.scala 44:32]
  wire [1:0] _T_1748; // @[LZD.scala 43:32]
  wire  _T_1749; // @[LZD.scala 39:14]
  wire  _T_1750; // @[LZD.scala 39:21]
  wire  _T_1751; // @[LZD.scala 39:30]
  wire  _T_1752; // @[LZD.scala 39:27]
  wire  _T_1753; // @[LZD.scala 39:25]
  wire [1:0] _T_1754; // @[Cat.scala 29:58]
  wire [1:0] _T_1755; // @[LZD.scala 44:32]
  wire  _T_1756; // @[LZD.scala 39:14]
  wire  _T_1757; // @[LZD.scala 39:21]
  wire  _T_1758; // @[LZD.scala 39:30]
  wire  _T_1759; // @[LZD.scala 39:27]
  wire  _T_1760; // @[LZD.scala 39:25]
  wire [1:0] _T_1761; // @[Cat.scala 29:58]
  wire  _T_1762; // @[Shift.scala 12:21]
  wire  _T_1763; // @[Shift.scala 12:21]
  wire  _T_1764; // @[LZD.scala 49:16]
  wire  _T_1765; // @[LZD.scala 49:27]
  wire  _T_1766; // @[LZD.scala 49:25]
  wire  _T_1767; // @[LZD.scala 49:47]
  wire  _T_1768; // @[LZD.scala 49:59]
  wire  _T_1769; // @[LZD.scala 49:35]
  wire [2:0] _T_1771; // @[Cat.scala 29:58]
  wire  _T_1772; // @[Shift.scala 12:21]
  wire  _T_1773; // @[Shift.scala 12:21]
  wire  _T_1774; // @[LZD.scala 49:16]
  wire  _T_1775; // @[LZD.scala 49:27]
  wire  _T_1776; // @[LZD.scala 49:25]
  wire [1:0] _T_1777; // @[LZD.scala 49:47]
  wire [1:0] _T_1778; // @[LZD.scala 49:59]
  wire [1:0] _T_1779; // @[LZD.scala 49:35]
  wire [3:0] _T_1781; // @[Cat.scala 29:58]
  wire [7:0] _T_1782; // @[LZD.scala 44:32]
  wire [3:0] _T_1783; // @[LZD.scala 43:32]
  wire [1:0] _T_1784; // @[LZD.scala 43:32]
  wire  _T_1785; // @[LZD.scala 39:14]
  wire  _T_1786; // @[LZD.scala 39:21]
  wire  _T_1787; // @[LZD.scala 39:30]
  wire  _T_1788; // @[LZD.scala 39:27]
  wire  _T_1789; // @[LZD.scala 39:25]
  wire [1:0] _T_1790; // @[Cat.scala 29:58]
  wire [1:0] _T_1791; // @[LZD.scala 44:32]
  wire  _T_1792; // @[LZD.scala 39:14]
  wire  _T_1793; // @[LZD.scala 39:21]
  wire  _T_1794; // @[LZD.scala 39:30]
  wire  _T_1795; // @[LZD.scala 39:27]
  wire  _T_1796; // @[LZD.scala 39:25]
  wire [1:0] _T_1797; // @[Cat.scala 29:58]
  wire  _T_1798; // @[Shift.scala 12:21]
  wire  _T_1799; // @[Shift.scala 12:21]
  wire  _T_1800; // @[LZD.scala 49:16]
  wire  _T_1801; // @[LZD.scala 49:27]
  wire  _T_1802; // @[LZD.scala 49:25]
  wire  _T_1803; // @[LZD.scala 49:47]
  wire  _T_1804; // @[LZD.scala 49:59]
  wire  _T_1805; // @[LZD.scala 49:35]
  wire [2:0] _T_1807; // @[Cat.scala 29:58]
  wire [3:0] _T_1808; // @[LZD.scala 44:32]
  wire [1:0] _T_1809; // @[LZD.scala 43:32]
  wire  _T_1810; // @[LZD.scala 39:14]
  wire  _T_1811; // @[LZD.scala 39:21]
  wire  _T_1812; // @[LZD.scala 39:30]
  wire  _T_1813; // @[LZD.scala 39:27]
  wire  _T_1814; // @[LZD.scala 39:25]
  wire [1:0] _T_1815; // @[Cat.scala 29:58]
  wire [1:0] _T_1816; // @[LZD.scala 44:32]
  wire  _T_1817; // @[LZD.scala 39:14]
  wire  _T_1818; // @[LZD.scala 39:21]
  wire  _T_1819; // @[LZD.scala 39:30]
  wire  _T_1820; // @[LZD.scala 39:27]
  wire  _T_1821; // @[LZD.scala 39:25]
  wire [1:0] _T_1822; // @[Cat.scala 29:58]
  wire  _T_1823; // @[Shift.scala 12:21]
  wire  _T_1824; // @[Shift.scala 12:21]
  wire  _T_1825; // @[LZD.scala 49:16]
  wire  _T_1826; // @[LZD.scala 49:27]
  wire  _T_1827; // @[LZD.scala 49:25]
  wire  _T_1828; // @[LZD.scala 49:47]
  wire  _T_1829; // @[LZD.scala 49:59]
  wire  _T_1830; // @[LZD.scala 49:35]
  wire [2:0] _T_1832; // @[Cat.scala 29:58]
  wire  _T_1833; // @[Shift.scala 12:21]
  wire  _T_1834; // @[Shift.scala 12:21]
  wire  _T_1835; // @[LZD.scala 49:16]
  wire  _T_1836; // @[LZD.scala 49:27]
  wire  _T_1837; // @[LZD.scala 49:25]
  wire [1:0] _T_1838; // @[LZD.scala 49:47]
  wire [1:0] _T_1839; // @[LZD.scala 49:59]
  wire [1:0] _T_1840; // @[LZD.scala 49:35]
  wire [3:0] _T_1842; // @[Cat.scala 29:58]
  wire  _T_1843; // @[Shift.scala 12:21]
  wire  _T_1844; // @[Shift.scala 12:21]
  wire  _T_1845; // @[LZD.scala 49:16]
  wire  _T_1846; // @[LZD.scala 49:27]
  wire  _T_1847; // @[LZD.scala 49:25]
  wire [2:0] _T_1848; // @[LZD.scala 49:47]
  wire [2:0] _T_1849; // @[LZD.scala 49:59]
  wire [2:0] _T_1850; // @[LZD.scala 49:35]
  wire [4:0] _T_1852; // @[Cat.scala 29:58]
  wire [15:0] _T_1853; // @[LZD.scala 44:32]
  wire [7:0] _T_1854; // @[LZD.scala 43:32]
  wire [3:0] _T_1855; // @[LZD.scala 43:32]
  wire [1:0] _T_1856; // @[LZD.scala 43:32]
  wire  _T_1857; // @[LZD.scala 39:14]
  wire  _T_1858; // @[LZD.scala 39:21]
  wire  _T_1859; // @[LZD.scala 39:30]
  wire  _T_1860; // @[LZD.scala 39:27]
  wire  _T_1861; // @[LZD.scala 39:25]
  wire [1:0] _T_1862; // @[Cat.scala 29:58]
  wire [1:0] _T_1863; // @[LZD.scala 44:32]
  wire  _T_1864; // @[LZD.scala 39:14]
  wire  _T_1865; // @[LZD.scala 39:21]
  wire  _T_1866; // @[LZD.scala 39:30]
  wire  _T_1867; // @[LZD.scala 39:27]
  wire  _T_1868; // @[LZD.scala 39:25]
  wire [1:0] _T_1869; // @[Cat.scala 29:58]
  wire  _T_1870; // @[Shift.scala 12:21]
  wire  _T_1871; // @[Shift.scala 12:21]
  wire  _T_1872; // @[LZD.scala 49:16]
  wire  _T_1873; // @[LZD.scala 49:27]
  wire  _T_1874; // @[LZD.scala 49:25]
  wire  _T_1875; // @[LZD.scala 49:47]
  wire  _T_1876; // @[LZD.scala 49:59]
  wire  _T_1877; // @[LZD.scala 49:35]
  wire [2:0] _T_1879; // @[Cat.scala 29:58]
  wire [3:0] _T_1880; // @[LZD.scala 44:32]
  wire [1:0] _T_1881; // @[LZD.scala 43:32]
  wire  _T_1882; // @[LZD.scala 39:14]
  wire  _T_1883; // @[LZD.scala 39:21]
  wire  _T_1884; // @[LZD.scala 39:30]
  wire  _T_1885; // @[LZD.scala 39:27]
  wire  _T_1886; // @[LZD.scala 39:25]
  wire [1:0] _T_1887; // @[Cat.scala 29:58]
  wire [1:0] _T_1888; // @[LZD.scala 44:32]
  wire  _T_1889; // @[LZD.scala 39:14]
  wire  _T_1890; // @[LZD.scala 39:21]
  wire  _T_1891; // @[LZD.scala 39:30]
  wire  _T_1892; // @[LZD.scala 39:27]
  wire  _T_1893; // @[LZD.scala 39:25]
  wire [1:0] _T_1894; // @[Cat.scala 29:58]
  wire  _T_1895; // @[Shift.scala 12:21]
  wire  _T_1896; // @[Shift.scala 12:21]
  wire  _T_1897; // @[LZD.scala 49:16]
  wire  _T_1898; // @[LZD.scala 49:27]
  wire  _T_1899; // @[LZD.scala 49:25]
  wire  _T_1900; // @[LZD.scala 49:47]
  wire  _T_1901; // @[LZD.scala 49:59]
  wire  _T_1902; // @[LZD.scala 49:35]
  wire [2:0] _T_1904; // @[Cat.scala 29:58]
  wire  _T_1905; // @[Shift.scala 12:21]
  wire  _T_1906; // @[Shift.scala 12:21]
  wire  _T_1907; // @[LZD.scala 49:16]
  wire  _T_1908; // @[LZD.scala 49:27]
  wire  _T_1909; // @[LZD.scala 49:25]
  wire [1:0] _T_1910; // @[LZD.scala 49:47]
  wire [1:0] _T_1911; // @[LZD.scala 49:59]
  wire [1:0] _T_1912; // @[LZD.scala 49:35]
  wire [3:0] _T_1914; // @[Cat.scala 29:58]
  wire [7:0] _T_1915; // @[LZD.scala 44:32]
  wire [3:0] _T_1916; // @[LZD.scala 43:32]
  wire [1:0] _T_1917; // @[LZD.scala 43:32]
  wire  _T_1918; // @[LZD.scala 39:14]
  wire  _T_1919; // @[LZD.scala 39:21]
  wire  _T_1920; // @[LZD.scala 39:30]
  wire  _T_1921; // @[LZD.scala 39:27]
  wire  _T_1922; // @[LZD.scala 39:25]
  wire [1:0] _T_1923; // @[Cat.scala 29:58]
  wire [1:0] _T_1924; // @[LZD.scala 44:32]
  wire  _T_1925; // @[LZD.scala 39:14]
  wire  _T_1926; // @[LZD.scala 39:21]
  wire  _T_1927; // @[LZD.scala 39:30]
  wire  _T_1928; // @[LZD.scala 39:27]
  wire  _T_1929; // @[LZD.scala 39:25]
  wire [1:0] _T_1930; // @[Cat.scala 29:58]
  wire  _T_1931; // @[Shift.scala 12:21]
  wire  _T_1932; // @[Shift.scala 12:21]
  wire  _T_1933; // @[LZD.scala 49:16]
  wire  _T_1934; // @[LZD.scala 49:27]
  wire  _T_1935; // @[LZD.scala 49:25]
  wire  _T_1936; // @[LZD.scala 49:47]
  wire  _T_1937; // @[LZD.scala 49:59]
  wire  _T_1938; // @[LZD.scala 49:35]
  wire [2:0] _T_1940; // @[Cat.scala 29:58]
  wire [3:0] _T_1941; // @[LZD.scala 44:32]
  wire [1:0] _T_1942; // @[LZD.scala 43:32]
  wire  _T_1943; // @[LZD.scala 39:14]
  wire  _T_1944; // @[LZD.scala 39:21]
  wire  _T_1945; // @[LZD.scala 39:30]
  wire  _T_1946; // @[LZD.scala 39:27]
  wire  _T_1947; // @[LZD.scala 39:25]
  wire [1:0] _T_1948; // @[Cat.scala 29:58]
  wire [1:0] _T_1949; // @[LZD.scala 44:32]
  wire  _T_1950; // @[LZD.scala 39:14]
  wire  _T_1951; // @[LZD.scala 39:21]
  wire  _T_1952; // @[LZD.scala 39:30]
  wire  _T_1953; // @[LZD.scala 39:27]
  wire  _T_1954; // @[LZD.scala 39:25]
  wire [1:0] _T_1955; // @[Cat.scala 29:58]
  wire  _T_1956; // @[Shift.scala 12:21]
  wire  _T_1957; // @[Shift.scala 12:21]
  wire  _T_1958; // @[LZD.scala 49:16]
  wire  _T_1959; // @[LZD.scala 49:27]
  wire  _T_1960; // @[LZD.scala 49:25]
  wire  _T_1961; // @[LZD.scala 49:47]
  wire  _T_1962; // @[LZD.scala 49:59]
  wire  _T_1963; // @[LZD.scala 49:35]
  wire [2:0] _T_1965; // @[Cat.scala 29:58]
  wire  _T_1966; // @[Shift.scala 12:21]
  wire  _T_1967; // @[Shift.scala 12:21]
  wire  _T_1968; // @[LZD.scala 49:16]
  wire  _T_1969; // @[LZD.scala 49:27]
  wire  _T_1970; // @[LZD.scala 49:25]
  wire [1:0] _T_1971; // @[LZD.scala 49:47]
  wire [1:0] _T_1972; // @[LZD.scala 49:59]
  wire [1:0] _T_1973; // @[LZD.scala 49:35]
  wire [3:0] _T_1975; // @[Cat.scala 29:58]
  wire  _T_1976; // @[Shift.scala 12:21]
  wire  _T_1977; // @[Shift.scala 12:21]
  wire  _T_1978; // @[LZD.scala 49:16]
  wire  _T_1979; // @[LZD.scala 49:27]
  wire  _T_1980; // @[LZD.scala 49:25]
  wire [2:0] _T_1981; // @[LZD.scala 49:47]
  wire [2:0] _T_1982; // @[LZD.scala 49:59]
  wire [2:0] _T_1983; // @[LZD.scala 49:35]
  wire [4:0] _T_1985; // @[Cat.scala 29:58]
  wire  _T_1986; // @[Shift.scala 12:21]
  wire  _T_1987; // @[Shift.scala 12:21]
  wire  _T_1988; // @[LZD.scala 49:16]
  wire  _T_1989; // @[LZD.scala 49:27]
  wire  _T_1990; // @[LZD.scala 49:25]
  wire [3:0] _T_1991; // @[LZD.scala 49:47]
  wire [3:0] _T_1992; // @[LZD.scala 49:59]
  wire [3:0] _T_1993; // @[LZD.scala 49:35]
  wire [5:0] _T_1995; // @[Cat.scala 29:58]
  wire [31:0] _T_1996; // @[LZD.scala 44:32]
  wire [15:0] _T_1997; // @[LZD.scala 43:32]
  wire [7:0] _T_1998; // @[LZD.scala 43:32]
  wire [3:0] _T_1999; // @[LZD.scala 43:32]
  wire [1:0] _T_2000; // @[LZD.scala 43:32]
  wire  _T_2001; // @[LZD.scala 39:14]
  wire  _T_2002; // @[LZD.scala 39:21]
  wire  _T_2003; // @[LZD.scala 39:30]
  wire  _T_2004; // @[LZD.scala 39:27]
  wire  _T_2005; // @[LZD.scala 39:25]
  wire [1:0] _T_2006; // @[Cat.scala 29:58]
  wire [1:0] _T_2007; // @[LZD.scala 44:32]
  wire  _T_2008; // @[LZD.scala 39:14]
  wire  _T_2009; // @[LZD.scala 39:21]
  wire  _T_2010; // @[LZD.scala 39:30]
  wire  _T_2011; // @[LZD.scala 39:27]
  wire  _T_2012; // @[LZD.scala 39:25]
  wire [1:0] _T_2013; // @[Cat.scala 29:58]
  wire  _T_2014; // @[Shift.scala 12:21]
  wire  _T_2015; // @[Shift.scala 12:21]
  wire  _T_2016; // @[LZD.scala 49:16]
  wire  _T_2017; // @[LZD.scala 49:27]
  wire  _T_2018; // @[LZD.scala 49:25]
  wire  _T_2019; // @[LZD.scala 49:47]
  wire  _T_2020; // @[LZD.scala 49:59]
  wire  _T_2021; // @[LZD.scala 49:35]
  wire [2:0] _T_2023; // @[Cat.scala 29:58]
  wire [3:0] _T_2024; // @[LZD.scala 44:32]
  wire [1:0] _T_2025; // @[LZD.scala 43:32]
  wire  _T_2026; // @[LZD.scala 39:14]
  wire  _T_2027; // @[LZD.scala 39:21]
  wire  _T_2028; // @[LZD.scala 39:30]
  wire  _T_2029; // @[LZD.scala 39:27]
  wire  _T_2030; // @[LZD.scala 39:25]
  wire [1:0] _T_2031; // @[Cat.scala 29:58]
  wire [1:0] _T_2032; // @[LZD.scala 44:32]
  wire  _T_2033; // @[LZD.scala 39:14]
  wire  _T_2034; // @[LZD.scala 39:21]
  wire  _T_2035; // @[LZD.scala 39:30]
  wire  _T_2036; // @[LZD.scala 39:27]
  wire  _T_2037; // @[LZD.scala 39:25]
  wire [1:0] _T_2038; // @[Cat.scala 29:58]
  wire  _T_2039; // @[Shift.scala 12:21]
  wire  _T_2040; // @[Shift.scala 12:21]
  wire  _T_2041; // @[LZD.scala 49:16]
  wire  _T_2042; // @[LZD.scala 49:27]
  wire  _T_2043; // @[LZD.scala 49:25]
  wire  _T_2044; // @[LZD.scala 49:47]
  wire  _T_2045; // @[LZD.scala 49:59]
  wire  _T_2046; // @[LZD.scala 49:35]
  wire [2:0] _T_2048; // @[Cat.scala 29:58]
  wire  _T_2049; // @[Shift.scala 12:21]
  wire  _T_2050; // @[Shift.scala 12:21]
  wire  _T_2051; // @[LZD.scala 49:16]
  wire  _T_2052; // @[LZD.scala 49:27]
  wire  _T_2053; // @[LZD.scala 49:25]
  wire [1:0] _T_2054; // @[LZD.scala 49:47]
  wire [1:0] _T_2055; // @[LZD.scala 49:59]
  wire [1:0] _T_2056; // @[LZD.scala 49:35]
  wire [3:0] _T_2058; // @[Cat.scala 29:58]
  wire [7:0] _T_2059; // @[LZD.scala 44:32]
  wire [3:0] _T_2060; // @[LZD.scala 43:32]
  wire [1:0] _T_2061; // @[LZD.scala 43:32]
  wire  _T_2062; // @[LZD.scala 39:14]
  wire  _T_2063; // @[LZD.scala 39:21]
  wire  _T_2064; // @[LZD.scala 39:30]
  wire  _T_2065; // @[LZD.scala 39:27]
  wire  _T_2066; // @[LZD.scala 39:25]
  wire [1:0] _T_2067; // @[Cat.scala 29:58]
  wire [1:0] _T_2068; // @[LZD.scala 44:32]
  wire  _T_2069; // @[LZD.scala 39:14]
  wire  _T_2070; // @[LZD.scala 39:21]
  wire  _T_2071; // @[LZD.scala 39:30]
  wire  _T_2072; // @[LZD.scala 39:27]
  wire  _T_2073; // @[LZD.scala 39:25]
  wire [1:0] _T_2074; // @[Cat.scala 29:58]
  wire  _T_2075; // @[Shift.scala 12:21]
  wire  _T_2076; // @[Shift.scala 12:21]
  wire  _T_2077; // @[LZD.scala 49:16]
  wire  _T_2078; // @[LZD.scala 49:27]
  wire  _T_2079; // @[LZD.scala 49:25]
  wire  _T_2080; // @[LZD.scala 49:47]
  wire  _T_2081; // @[LZD.scala 49:59]
  wire  _T_2082; // @[LZD.scala 49:35]
  wire [2:0] _T_2084; // @[Cat.scala 29:58]
  wire [3:0] _T_2085; // @[LZD.scala 44:32]
  wire [1:0] _T_2086; // @[LZD.scala 43:32]
  wire  _T_2087; // @[LZD.scala 39:14]
  wire  _T_2088; // @[LZD.scala 39:21]
  wire  _T_2089; // @[LZD.scala 39:30]
  wire  _T_2090; // @[LZD.scala 39:27]
  wire  _T_2091; // @[LZD.scala 39:25]
  wire [1:0] _T_2092; // @[Cat.scala 29:58]
  wire [1:0] _T_2093; // @[LZD.scala 44:32]
  wire  _T_2094; // @[LZD.scala 39:14]
  wire  _T_2095; // @[LZD.scala 39:21]
  wire  _T_2096; // @[LZD.scala 39:30]
  wire  _T_2097; // @[LZD.scala 39:27]
  wire  _T_2098; // @[LZD.scala 39:25]
  wire [1:0] _T_2099; // @[Cat.scala 29:58]
  wire  _T_2100; // @[Shift.scala 12:21]
  wire  _T_2101; // @[Shift.scala 12:21]
  wire  _T_2102; // @[LZD.scala 49:16]
  wire  _T_2103; // @[LZD.scala 49:27]
  wire  _T_2104; // @[LZD.scala 49:25]
  wire  _T_2105; // @[LZD.scala 49:47]
  wire  _T_2106; // @[LZD.scala 49:59]
  wire  _T_2107; // @[LZD.scala 49:35]
  wire [2:0] _T_2109; // @[Cat.scala 29:58]
  wire  _T_2110; // @[Shift.scala 12:21]
  wire  _T_2111; // @[Shift.scala 12:21]
  wire  _T_2112; // @[LZD.scala 49:16]
  wire  _T_2113; // @[LZD.scala 49:27]
  wire  _T_2114; // @[LZD.scala 49:25]
  wire [1:0] _T_2115; // @[LZD.scala 49:47]
  wire [1:0] _T_2116; // @[LZD.scala 49:59]
  wire [1:0] _T_2117; // @[LZD.scala 49:35]
  wire [3:0] _T_2119; // @[Cat.scala 29:58]
  wire  _T_2120; // @[Shift.scala 12:21]
  wire  _T_2121; // @[Shift.scala 12:21]
  wire  _T_2122; // @[LZD.scala 49:16]
  wire  _T_2123; // @[LZD.scala 49:27]
  wire  _T_2124; // @[LZD.scala 49:25]
  wire [2:0] _T_2125; // @[LZD.scala 49:47]
  wire [2:0] _T_2126; // @[LZD.scala 49:59]
  wire [2:0] _T_2127; // @[LZD.scala 49:35]
  wire [4:0] _T_2129; // @[Cat.scala 29:58]
  wire [15:0] _T_2130; // @[LZD.scala 44:32]
  wire [7:0] _T_2131; // @[LZD.scala 43:32]
  wire [3:0] _T_2132; // @[LZD.scala 43:32]
  wire [1:0] _T_2133; // @[LZD.scala 43:32]
  wire  _T_2134; // @[LZD.scala 39:14]
  wire  _T_2135; // @[LZD.scala 39:21]
  wire  _T_2136; // @[LZD.scala 39:30]
  wire  _T_2137; // @[LZD.scala 39:27]
  wire  _T_2138; // @[LZD.scala 39:25]
  wire [1:0] _T_2139; // @[Cat.scala 29:58]
  wire [1:0] _T_2140; // @[LZD.scala 44:32]
  wire  _T_2141; // @[LZD.scala 39:14]
  wire  _T_2142; // @[LZD.scala 39:21]
  wire  _T_2143; // @[LZD.scala 39:30]
  wire  _T_2144; // @[LZD.scala 39:27]
  wire  _T_2145; // @[LZD.scala 39:25]
  wire [1:0] _T_2146; // @[Cat.scala 29:58]
  wire  _T_2147; // @[Shift.scala 12:21]
  wire  _T_2148; // @[Shift.scala 12:21]
  wire  _T_2149; // @[LZD.scala 49:16]
  wire  _T_2150; // @[LZD.scala 49:27]
  wire  _T_2151; // @[LZD.scala 49:25]
  wire  _T_2152; // @[LZD.scala 49:47]
  wire  _T_2153; // @[LZD.scala 49:59]
  wire  _T_2154; // @[LZD.scala 49:35]
  wire [2:0] _T_2156; // @[Cat.scala 29:58]
  wire [3:0] _T_2157; // @[LZD.scala 44:32]
  wire [1:0] _T_2158; // @[LZD.scala 43:32]
  wire  _T_2159; // @[LZD.scala 39:14]
  wire  _T_2160; // @[LZD.scala 39:21]
  wire  _T_2161; // @[LZD.scala 39:30]
  wire  _T_2162; // @[LZD.scala 39:27]
  wire  _T_2163; // @[LZD.scala 39:25]
  wire [1:0] _T_2164; // @[Cat.scala 29:58]
  wire [1:0] _T_2165; // @[LZD.scala 44:32]
  wire  _T_2166; // @[LZD.scala 39:14]
  wire  _T_2167; // @[LZD.scala 39:21]
  wire  _T_2168; // @[LZD.scala 39:30]
  wire  _T_2169; // @[LZD.scala 39:27]
  wire  _T_2170; // @[LZD.scala 39:25]
  wire [1:0] _T_2171; // @[Cat.scala 29:58]
  wire  _T_2172; // @[Shift.scala 12:21]
  wire  _T_2173; // @[Shift.scala 12:21]
  wire  _T_2174; // @[LZD.scala 49:16]
  wire  _T_2175; // @[LZD.scala 49:27]
  wire  _T_2176; // @[LZD.scala 49:25]
  wire  _T_2177; // @[LZD.scala 49:47]
  wire  _T_2178; // @[LZD.scala 49:59]
  wire  _T_2179; // @[LZD.scala 49:35]
  wire [2:0] _T_2181; // @[Cat.scala 29:58]
  wire  _T_2182; // @[Shift.scala 12:21]
  wire  _T_2183; // @[Shift.scala 12:21]
  wire  _T_2184; // @[LZD.scala 49:16]
  wire  _T_2185; // @[LZD.scala 49:27]
  wire  _T_2186; // @[LZD.scala 49:25]
  wire [1:0] _T_2187; // @[LZD.scala 49:47]
  wire [1:0] _T_2188; // @[LZD.scala 49:59]
  wire [1:0] _T_2189; // @[LZD.scala 49:35]
  wire [3:0] _T_2191; // @[Cat.scala 29:58]
  wire [7:0] _T_2192; // @[LZD.scala 44:32]
  wire [3:0] _T_2193; // @[LZD.scala 43:32]
  wire [1:0] _T_2194; // @[LZD.scala 43:32]
  wire  _T_2195; // @[LZD.scala 39:14]
  wire  _T_2196; // @[LZD.scala 39:21]
  wire  _T_2197; // @[LZD.scala 39:30]
  wire  _T_2198; // @[LZD.scala 39:27]
  wire  _T_2199; // @[LZD.scala 39:25]
  wire [1:0] _T_2200; // @[Cat.scala 29:58]
  wire [1:0] _T_2201; // @[LZD.scala 44:32]
  wire  _T_2202; // @[LZD.scala 39:14]
  wire  _T_2203; // @[LZD.scala 39:21]
  wire  _T_2204; // @[LZD.scala 39:30]
  wire  _T_2205; // @[LZD.scala 39:27]
  wire  _T_2206; // @[LZD.scala 39:25]
  wire [1:0] _T_2207; // @[Cat.scala 29:58]
  wire  _T_2208; // @[Shift.scala 12:21]
  wire  _T_2209; // @[Shift.scala 12:21]
  wire  _T_2210; // @[LZD.scala 49:16]
  wire  _T_2211; // @[LZD.scala 49:27]
  wire  _T_2212; // @[LZD.scala 49:25]
  wire  _T_2213; // @[LZD.scala 49:47]
  wire  _T_2214; // @[LZD.scala 49:59]
  wire  _T_2215; // @[LZD.scala 49:35]
  wire [2:0] _T_2217; // @[Cat.scala 29:58]
  wire [3:0] _T_2218; // @[LZD.scala 44:32]
  wire [1:0] _T_2219; // @[LZD.scala 43:32]
  wire  _T_2220; // @[LZD.scala 39:14]
  wire  _T_2221; // @[LZD.scala 39:21]
  wire  _T_2222; // @[LZD.scala 39:30]
  wire  _T_2223; // @[LZD.scala 39:27]
  wire  _T_2224; // @[LZD.scala 39:25]
  wire [1:0] _T_2225; // @[Cat.scala 29:58]
  wire [1:0] _T_2226; // @[LZD.scala 44:32]
  wire  _T_2227; // @[LZD.scala 39:14]
  wire  _T_2228; // @[LZD.scala 39:21]
  wire  _T_2229; // @[LZD.scala 39:30]
  wire  _T_2230; // @[LZD.scala 39:27]
  wire  _T_2231; // @[LZD.scala 39:25]
  wire [1:0] _T_2232; // @[Cat.scala 29:58]
  wire  _T_2233; // @[Shift.scala 12:21]
  wire  _T_2234; // @[Shift.scala 12:21]
  wire  _T_2235; // @[LZD.scala 49:16]
  wire  _T_2236; // @[LZD.scala 49:27]
  wire  _T_2237; // @[LZD.scala 49:25]
  wire  _T_2238; // @[LZD.scala 49:47]
  wire  _T_2239; // @[LZD.scala 49:59]
  wire  _T_2240; // @[LZD.scala 49:35]
  wire [2:0] _T_2242; // @[Cat.scala 29:58]
  wire  _T_2243; // @[Shift.scala 12:21]
  wire  _T_2244; // @[Shift.scala 12:21]
  wire  _T_2245; // @[LZD.scala 49:16]
  wire  _T_2246; // @[LZD.scala 49:27]
  wire  _T_2247; // @[LZD.scala 49:25]
  wire [1:0] _T_2248; // @[LZD.scala 49:47]
  wire [1:0] _T_2249; // @[LZD.scala 49:59]
  wire [1:0] _T_2250; // @[LZD.scala 49:35]
  wire [3:0] _T_2252; // @[Cat.scala 29:58]
  wire  _T_2253; // @[Shift.scala 12:21]
  wire  _T_2254; // @[Shift.scala 12:21]
  wire  _T_2255; // @[LZD.scala 49:16]
  wire  _T_2256; // @[LZD.scala 49:27]
  wire  _T_2257; // @[LZD.scala 49:25]
  wire [2:0] _T_2258; // @[LZD.scala 49:47]
  wire [2:0] _T_2259; // @[LZD.scala 49:59]
  wire [2:0] _T_2260; // @[LZD.scala 49:35]
  wire [4:0] _T_2262; // @[Cat.scala 29:58]
  wire  _T_2263; // @[Shift.scala 12:21]
  wire  _T_2264; // @[Shift.scala 12:21]
  wire  _T_2265; // @[LZD.scala 49:16]
  wire  _T_2266; // @[LZD.scala 49:27]
  wire  _T_2267; // @[LZD.scala 49:25]
  wire [3:0] _T_2268; // @[LZD.scala 49:47]
  wire [3:0] _T_2269; // @[LZD.scala 49:59]
  wire [3:0] _T_2270; // @[LZD.scala 49:35]
  wire [5:0] _T_2272; // @[Cat.scala 29:58]
  wire  _T_2273; // @[Shift.scala 12:21]
  wire  _T_2274; // @[Shift.scala 12:21]
  wire  _T_2275; // @[LZD.scala 49:16]
  wire  _T_2276; // @[LZD.scala 49:27]
  wire  _T_2277; // @[LZD.scala 49:25]
  wire [4:0] _T_2278; // @[LZD.scala 49:47]
  wire [4:0] _T_2279; // @[LZD.scala 49:59]
  wire [4:0] _T_2280; // @[LZD.scala 49:35]
  wire [6:0] _T_2282; // @[Cat.scala 29:58]
  wire  _T_2283; // @[Shift.scala 12:21]
  wire  _T_2284; // @[Shift.scala 12:21]
  wire  _T_2285; // @[LZD.scala 49:16]
  wire  _T_2286; // @[LZD.scala 49:27]
  wire  _T_2287; // @[LZD.scala 49:25]
  wire [5:0] _T_2288; // @[LZD.scala 49:47]
  wire [5:0] _T_2289; // @[LZD.scala 49:59]
  wire [5:0] _T_2290; // @[LZD.scala 49:35]
  wire [7:0] _T_2292; // @[Cat.scala 29:58]
  wire  _T_2293; // @[Shift.scala 12:21]
  wire  _T_2294; // @[Shift.scala 12:21]
  wire  _T_2295; // @[LZD.scala 49:16]
  wire  _T_2296; // @[LZD.scala 49:27]
  wire  _T_2297; // @[LZD.scala 49:25]
  wire [6:0] _T_2298; // @[LZD.scala 49:47]
  wire [6:0] _T_2299; // @[LZD.scala 49:59]
  wire [6:0] _T_2300; // @[LZD.scala 49:35]
  wire [8:0] _T_2302; // @[Cat.scala 29:58]
  wire [56:0] _T_2303; // @[LZD.scala 44:32]
  wire [31:0] _T_2304; // @[LZD.scala 43:32]
  wire [15:0] _T_2305; // @[LZD.scala 43:32]
  wire [7:0] _T_2306; // @[LZD.scala 43:32]
  wire [3:0] _T_2307; // @[LZD.scala 43:32]
  wire [1:0] _T_2308; // @[LZD.scala 43:32]
  wire  _T_2309; // @[LZD.scala 39:14]
  wire  _T_2310; // @[LZD.scala 39:21]
  wire  _T_2311; // @[LZD.scala 39:30]
  wire  _T_2312; // @[LZD.scala 39:27]
  wire  _T_2313; // @[LZD.scala 39:25]
  wire [1:0] _T_2314; // @[Cat.scala 29:58]
  wire [1:0] _T_2315; // @[LZD.scala 44:32]
  wire  _T_2316; // @[LZD.scala 39:14]
  wire  _T_2317; // @[LZD.scala 39:21]
  wire  _T_2318; // @[LZD.scala 39:30]
  wire  _T_2319; // @[LZD.scala 39:27]
  wire  _T_2320; // @[LZD.scala 39:25]
  wire [1:0] _T_2321; // @[Cat.scala 29:58]
  wire  _T_2322; // @[Shift.scala 12:21]
  wire  _T_2323; // @[Shift.scala 12:21]
  wire  _T_2324; // @[LZD.scala 49:16]
  wire  _T_2325; // @[LZD.scala 49:27]
  wire  _T_2326; // @[LZD.scala 49:25]
  wire  _T_2327; // @[LZD.scala 49:47]
  wire  _T_2328; // @[LZD.scala 49:59]
  wire  _T_2329; // @[LZD.scala 49:35]
  wire [2:0] _T_2331; // @[Cat.scala 29:58]
  wire [3:0] _T_2332; // @[LZD.scala 44:32]
  wire [1:0] _T_2333; // @[LZD.scala 43:32]
  wire  _T_2334; // @[LZD.scala 39:14]
  wire  _T_2335; // @[LZD.scala 39:21]
  wire  _T_2336; // @[LZD.scala 39:30]
  wire  _T_2337; // @[LZD.scala 39:27]
  wire  _T_2338; // @[LZD.scala 39:25]
  wire [1:0] _T_2339; // @[Cat.scala 29:58]
  wire [1:0] _T_2340; // @[LZD.scala 44:32]
  wire  _T_2341; // @[LZD.scala 39:14]
  wire  _T_2342; // @[LZD.scala 39:21]
  wire  _T_2343; // @[LZD.scala 39:30]
  wire  _T_2344; // @[LZD.scala 39:27]
  wire  _T_2345; // @[LZD.scala 39:25]
  wire [1:0] _T_2346; // @[Cat.scala 29:58]
  wire  _T_2347; // @[Shift.scala 12:21]
  wire  _T_2348; // @[Shift.scala 12:21]
  wire  _T_2349; // @[LZD.scala 49:16]
  wire  _T_2350; // @[LZD.scala 49:27]
  wire  _T_2351; // @[LZD.scala 49:25]
  wire  _T_2352; // @[LZD.scala 49:47]
  wire  _T_2353; // @[LZD.scala 49:59]
  wire  _T_2354; // @[LZD.scala 49:35]
  wire [2:0] _T_2356; // @[Cat.scala 29:58]
  wire  _T_2357; // @[Shift.scala 12:21]
  wire  _T_2358; // @[Shift.scala 12:21]
  wire  _T_2359; // @[LZD.scala 49:16]
  wire  _T_2360; // @[LZD.scala 49:27]
  wire  _T_2361; // @[LZD.scala 49:25]
  wire [1:0] _T_2362; // @[LZD.scala 49:47]
  wire [1:0] _T_2363; // @[LZD.scala 49:59]
  wire [1:0] _T_2364; // @[LZD.scala 49:35]
  wire [3:0] _T_2366; // @[Cat.scala 29:58]
  wire [7:0] _T_2367; // @[LZD.scala 44:32]
  wire [3:0] _T_2368; // @[LZD.scala 43:32]
  wire [1:0] _T_2369; // @[LZD.scala 43:32]
  wire  _T_2370; // @[LZD.scala 39:14]
  wire  _T_2371; // @[LZD.scala 39:21]
  wire  _T_2372; // @[LZD.scala 39:30]
  wire  _T_2373; // @[LZD.scala 39:27]
  wire  _T_2374; // @[LZD.scala 39:25]
  wire [1:0] _T_2375; // @[Cat.scala 29:58]
  wire [1:0] _T_2376; // @[LZD.scala 44:32]
  wire  _T_2377; // @[LZD.scala 39:14]
  wire  _T_2378; // @[LZD.scala 39:21]
  wire  _T_2379; // @[LZD.scala 39:30]
  wire  _T_2380; // @[LZD.scala 39:27]
  wire  _T_2381; // @[LZD.scala 39:25]
  wire [1:0] _T_2382; // @[Cat.scala 29:58]
  wire  _T_2383; // @[Shift.scala 12:21]
  wire  _T_2384; // @[Shift.scala 12:21]
  wire  _T_2385; // @[LZD.scala 49:16]
  wire  _T_2386; // @[LZD.scala 49:27]
  wire  _T_2387; // @[LZD.scala 49:25]
  wire  _T_2388; // @[LZD.scala 49:47]
  wire  _T_2389; // @[LZD.scala 49:59]
  wire  _T_2390; // @[LZD.scala 49:35]
  wire [2:0] _T_2392; // @[Cat.scala 29:58]
  wire [3:0] _T_2393; // @[LZD.scala 44:32]
  wire [1:0] _T_2394; // @[LZD.scala 43:32]
  wire  _T_2395; // @[LZD.scala 39:14]
  wire  _T_2396; // @[LZD.scala 39:21]
  wire  _T_2397; // @[LZD.scala 39:30]
  wire  _T_2398; // @[LZD.scala 39:27]
  wire  _T_2399; // @[LZD.scala 39:25]
  wire [1:0] _T_2400; // @[Cat.scala 29:58]
  wire [1:0] _T_2401; // @[LZD.scala 44:32]
  wire  _T_2402; // @[LZD.scala 39:14]
  wire  _T_2403; // @[LZD.scala 39:21]
  wire  _T_2404; // @[LZD.scala 39:30]
  wire  _T_2405; // @[LZD.scala 39:27]
  wire  _T_2406; // @[LZD.scala 39:25]
  wire [1:0] _T_2407; // @[Cat.scala 29:58]
  wire  _T_2408; // @[Shift.scala 12:21]
  wire  _T_2409; // @[Shift.scala 12:21]
  wire  _T_2410; // @[LZD.scala 49:16]
  wire  _T_2411; // @[LZD.scala 49:27]
  wire  _T_2412; // @[LZD.scala 49:25]
  wire  _T_2413; // @[LZD.scala 49:47]
  wire  _T_2414; // @[LZD.scala 49:59]
  wire  _T_2415; // @[LZD.scala 49:35]
  wire [2:0] _T_2417; // @[Cat.scala 29:58]
  wire  _T_2418; // @[Shift.scala 12:21]
  wire  _T_2419; // @[Shift.scala 12:21]
  wire  _T_2420; // @[LZD.scala 49:16]
  wire  _T_2421; // @[LZD.scala 49:27]
  wire  _T_2422; // @[LZD.scala 49:25]
  wire [1:0] _T_2423; // @[LZD.scala 49:47]
  wire [1:0] _T_2424; // @[LZD.scala 49:59]
  wire [1:0] _T_2425; // @[LZD.scala 49:35]
  wire [3:0] _T_2427; // @[Cat.scala 29:58]
  wire  _T_2428; // @[Shift.scala 12:21]
  wire  _T_2429; // @[Shift.scala 12:21]
  wire  _T_2430; // @[LZD.scala 49:16]
  wire  _T_2431; // @[LZD.scala 49:27]
  wire  _T_2432; // @[LZD.scala 49:25]
  wire [2:0] _T_2433; // @[LZD.scala 49:47]
  wire [2:0] _T_2434; // @[LZD.scala 49:59]
  wire [2:0] _T_2435; // @[LZD.scala 49:35]
  wire [4:0] _T_2437; // @[Cat.scala 29:58]
  wire [15:0] _T_2438; // @[LZD.scala 44:32]
  wire [7:0] _T_2439; // @[LZD.scala 43:32]
  wire [3:0] _T_2440; // @[LZD.scala 43:32]
  wire [1:0] _T_2441; // @[LZD.scala 43:32]
  wire  _T_2442; // @[LZD.scala 39:14]
  wire  _T_2443; // @[LZD.scala 39:21]
  wire  _T_2444; // @[LZD.scala 39:30]
  wire  _T_2445; // @[LZD.scala 39:27]
  wire  _T_2446; // @[LZD.scala 39:25]
  wire [1:0] _T_2447; // @[Cat.scala 29:58]
  wire [1:0] _T_2448; // @[LZD.scala 44:32]
  wire  _T_2449; // @[LZD.scala 39:14]
  wire  _T_2450; // @[LZD.scala 39:21]
  wire  _T_2451; // @[LZD.scala 39:30]
  wire  _T_2452; // @[LZD.scala 39:27]
  wire  _T_2453; // @[LZD.scala 39:25]
  wire [1:0] _T_2454; // @[Cat.scala 29:58]
  wire  _T_2455; // @[Shift.scala 12:21]
  wire  _T_2456; // @[Shift.scala 12:21]
  wire  _T_2457; // @[LZD.scala 49:16]
  wire  _T_2458; // @[LZD.scala 49:27]
  wire  _T_2459; // @[LZD.scala 49:25]
  wire  _T_2460; // @[LZD.scala 49:47]
  wire  _T_2461; // @[LZD.scala 49:59]
  wire  _T_2462; // @[LZD.scala 49:35]
  wire [2:0] _T_2464; // @[Cat.scala 29:58]
  wire [3:0] _T_2465; // @[LZD.scala 44:32]
  wire [1:0] _T_2466; // @[LZD.scala 43:32]
  wire  _T_2467; // @[LZD.scala 39:14]
  wire  _T_2468; // @[LZD.scala 39:21]
  wire  _T_2469; // @[LZD.scala 39:30]
  wire  _T_2470; // @[LZD.scala 39:27]
  wire  _T_2471; // @[LZD.scala 39:25]
  wire [1:0] _T_2472; // @[Cat.scala 29:58]
  wire [1:0] _T_2473; // @[LZD.scala 44:32]
  wire  _T_2474; // @[LZD.scala 39:14]
  wire  _T_2475; // @[LZD.scala 39:21]
  wire  _T_2476; // @[LZD.scala 39:30]
  wire  _T_2477; // @[LZD.scala 39:27]
  wire  _T_2478; // @[LZD.scala 39:25]
  wire [1:0] _T_2479; // @[Cat.scala 29:58]
  wire  _T_2480; // @[Shift.scala 12:21]
  wire  _T_2481; // @[Shift.scala 12:21]
  wire  _T_2482; // @[LZD.scala 49:16]
  wire  _T_2483; // @[LZD.scala 49:27]
  wire  _T_2484; // @[LZD.scala 49:25]
  wire  _T_2485; // @[LZD.scala 49:47]
  wire  _T_2486; // @[LZD.scala 49:59]
  wire  _T_2487; // @[LZD.scala 49:35]
  wire [2:0] _T_2489; // @[Cat.scala 29:58]
  wire  _T_2490; // @[Shift.scala 12:21]
  wire  _T_2491; // @[Shift.scala 12:21]
  wire  _T_2492; // @[LZD.scala 49:16]
  wire  _T_2493; // @[LZD.scala 49:27]
  wire  _T_2494; // @[LZD.scala 49:25]
  wire [1:0] _T_2495; // @[LZD.scala 49:47]
  wire [1:0] _T_2496; // @[LZD.scala 49:59]
  wire [1:0] _T_2497; // @[LZD.scala 49:35]
  wire [3:0] _T_2499; // @[Cat.scala 29:58]
  wire [7:0] _T_2500; // @[LZD.scala 44:32]
  wire [3:0] _T_2501; // @[LZD.scala 43:32]
  wire [1:0] _T_2502; // @[LZD.scala 43:32]
  wire  _T_2503; // @[LZD.scala 39:14]
  wire  _T_2504; // @[LZD.scala 39:21]
  wire  _T_2505; // @[LZD.scala 39:30]
  wire  _T_2506; // @[LZD.scala 39:27]
  wire  _T_2507; // @[LZD.scala 39:25]
  wire [1:0] _T_2508; // @[Cat.scala 29:58]
  wire [1:0] _T_2509; // @[LZD.scala 44:32]
  wire  _T_2510; // @[LZD.scala 39:14]
  wire  _T_2511; // @[LZD.scala 39:21]
  wire  _T_2512; // @[LZD.scala 39:30]
  wire  _T_2513; // @[LZD.scala 39:27]
  wire  _T_2514; // @[LZD.scala 39:25]
  wire [1:0] _T_2515; // @[Cat.scala 29:58]
  wire  _T_2516; // @[Shift.scala 12:21]
  wire  _T_2517; // @[Shift.scala 12:21]
  wire  _T_2518; // @[LZD.scala 49:16]
  wire  _T_2519; // @[LZD.scala 49:27]
  wire  _T_2520; // @[LZD.scala 49:25]
  wire  _T_2521; // @[LZD.scala 49:47]
  wire  _T_2522; // @[LZD.scala 49:59]
  wire  _T_2523; // @[LZD.scala 49:35]
  wire [2:0] _T_2525; // @[Cat.scala 29:58]
  wire [3:0] _T_2526; // @[LZD.scala 44:32]
  wire [1:0] _T_2527; // @[LZD.scala 43:32]
  wire  _T_2528; // @[LZD.scala 39:14]
  wire  _T_2529; // @[LZD.scala 39:21]
  wire  _T_2530; // @[LZD.scala 39:30]
  wire  _T_2531; // @[LZD.scala 39:27]
  wire  _T_2532; // @[LZD.scala 39:25]
  wire [1:0] _T_2533; // @[Cat.scala 29:58]
  wire [1:0] _T_2534; // @[LZD.scala 44:32]
  wire  _T_2535; // @[LZD.scala 39:14]
  wire  _T_2536; // @[LZD.scala 39:21]
  wire  _T_2537; // @[LZD.scala 39:30]
  wire  _T_2538; // @[LZD.scala 39:27]
  wire  _T_2539; // @[LZD.scala 39:25]
  wire [1:0] _T_2540; // @[Cat.scala 29:58]
  wire  _T_2541; // @[Shift.scala 12:21]
  wire  _T_2542; // @[Shift.scala 12:21]
  wire  _T_2543; // @[LZD.scala 49:16]
  wire  _T_2544; // @[LZD.scala 49:27]
  wire  _T_2545; // @[LZD.scala 49:25]
  wire  _T_2546; // @[LZD.scala 49:47]
  wire  _T_2547; // @[LZD.scala 49:59]
  wire  _T_2548; // @[LZD.scala 49:35]
  wire [2:0] _T_2550; // @[Cat.scala 29:58]
  wire  _T_2551; // @[Shift.scala 12:21]
  wire  _T_2552; // @[Shift.scala 12:21]
  wire  _T_2553; // @[LZD.scala 49:16]
  wire  _T_2554; // @[LZD.scala 49:27]
  wire  _T_2555; // @[LZD.scala 49:25]
  wire [1:0] _T_2556; // @[LZD.scala 49:47]
  wire [1:0] _T_2557; // @[LZD.scala 49:59]
  wire [1:0] _T_2558; // @[LZD.scala 49:35]
  wire [3:0] _T_2560; // @[Cat.scala 29:58]
  wire  _T_2561; // @[Shift.scala 12:21]
  wire  _T_2562; // @[Shift.scala 12:21]
  wire  _T_2563; // @[LZD.scala 49:16]
  wire  _T_2564; // @[LZD.scala 49:27]
  wire  _T_2565; // @[LZD.scala 49:25]
  wire [2:0] _T_2566; // @[LZD.scala 49:47]
  wire [2:0] _T_2567; // @[LZD.scala 49:59]
  wire [2:0] _T_2568; // @[LZD.scala 49:35]
  wire [4:0] _T_2570; // @[Cat.scala 29:58]
  wire  _T_2571; // @[Shift.scala 12:21]
  wire  _T_2572; // @[Shift.scala 12:21]
  wire  _T_2573; // @[LZD.scala 49:16]
  wire  _T_2574; // @[LZD.scala 49:27]
  wire  _T_2575; // @[LZD.scala 49:25]
  wire [3:0] _T_2576; // @[LZD.scala 49:47]
  wire [3:0] _T_2577; // @[LZD.scala 49:59]
  wire [3:0] _T_2578; // @[LZD.scala 49:35]
  wire [5:0] _T_2580; // @[Cat.scala 29:58]
  wire [24:0] _T_2581; // @[LZD.scala 44:32]
  wire [15:0] _T_2582; // @[LZD.scala 43:32]
  wire [7:0] _T_2583; // @[LZD.scala 43:32]
  wire [3:0] _T_2584; // @[LZD.scala 43:32]
  wire [1:0] _T_2585; // @[LZD.scala 43:32]
  wire  _T_2586; // @[LZD.scala 39:14]
  wire  _T_2587; // @[LZD.scala 39:21]
  wire  _T_2588; // @[LZD.scala 39:30]
  wire  _T_2589; // @[LZD.scala 39:27]
  wire  _T_2590; // @[LZD.scala 39:25]
  wire [1:0] _T_2591; // @[Cat.scala 29:58]
  wire [1:0] _T_2592; // @[LZD.scala 44:32]
  wire  _T_2593; // @[LZD.scala 39:14]
  wire  _T_2594; // @[LZD.scala 39:21]
  wire  _T_2595; // @[LZD.scala 39:30]
  wire  _T_2596; // @[LZD.scala 39:27]
  wire  _T_2597; // @[LZD.scala 39:25]
  wire [1:0] _T_2598; // @[Cat.scala 29:58]
  wire  _T_2599; // @[Shift.scala 12:21]
  wire  _T_2600; // @[Shift.scala 12:21]
  wire  _T_2601; // @[LZD.scala 49:16]
  wire  _T_2602; // @[LZD.scala 49:27]
  wire  _T_2603; // @[LZD.scala 49:25]
  wire  _T_2604; // @[LZD.scala 49:47]
  wire  _T_2605; // @[LZD.scala 49:59]
  wire  _T_2606; // @[LZD.scala 49:35]
  wire [2:0] _T_2608; // @[Cat.scala 29:58]
  wire [3:0] _T_2609; // @[LZD.scala 44:32]
  wire [1:0] _T_2610; // @[LZD.scala 43:32]
  wire  _T_2611; // @[LZD.scala 39:14]
  wire  _T_2612; // @[LZD.scala 39:21]
  wire  _T_2613; // @[LZD.scala 39:30]
  wire  _T_2614; // @[LZD.scala 39:27]
  wire  _T_2615; // @[LZD.scala 39:25]
  wire [1:0] _T_2616; // @[Cat.scala 29:58]
  wire [1:0] _T_2617; // @[LZD.scala 44:32]
  wire  _T_2618; // @[LZD.scala 39:14]
  wire  _T_2619; // @[LZD.scala 39:21]
  wire  _T_2620; // @[LZD.scala 39:30]
  wire  _T_2621; // @[LZD.scala 39:27]
  wire  _T_2622; // @[LZD.scala 39:25]
  wire [1:0] _T_2623; // @[Cat.scala 29:58]
  wire  _T_2624; // @[Shift.scala 12:21]
  wire  _T_2625; // @[Shift.scala 12:21]
  wire  _T_2626; // @[LZD.scala 49:16]
  wire  _T_2627; // @[LZD.scala 49:27]
  wire  _T_2628; // @[LZD.scala 49:25]
  wire  _T_2629; // @[LZD.scala 49:47]
  wire  _T_2630; // @[LZD.scala 49:59]
  wire  _T_2631; // @[LZD.scala 49:35]
  wire [2:0] _T_2633; // @[Cat.scala 29:58]
  wire  _T_2634; // @[Shift.scala 12:21]
  wire  _T_2635; // @[Shift.scala 12:21]
  wire  _T_2636; // @[LZD.scala 49:16]
  wire  _T_2637; // @[LZD.scala 49:27]
  wire  _T_2638; // @[LZD.scala 49:25]
  wire [1:0] _T_2639; // @[LZD.scala 49:47]
  wire [1:0] _T_2640; // @[LZD.scala 49:59]
  wire [1:0] _T_2641; // @[LZD.scala 49:35]
  wire [3:0] _T_2643; // @[Cat.scala 29:58]
  wire [7:0] _T_2644; // @[LZD.scala 44:32]
  wire [3:0] _T_2645; // @[LZD.scala 43:32]
  wire [1:0] _T_2646; // @[LZD.scala 43:32]
  wire  _T_2647; // @[LZD.scala 39:14]
  wire  _T_2648; // @[LZD.scala 39:21]
  wire  _T_2649; // @[LZD.scala 39:30]
  wire  _T_2650; // @[LZD.scala 39:27]
  wire  _T_2651; // @[LZD.scala 39:25]
  wire [1:0] _T_2652; // @[Cat.scala 29:58]
  wire [1:0] _T_2653; // @[LZD.scala 44:32]
  wire  _T_2654; // @[LZD.scala 39:14]
  wire  _T_2655; // @[LZD.scala 39:21]
  wire  _T_2656; // @[LZD.scala 39:30]
  wire  _T_2657; // @[LZD.scala 39:27]
  wire  _T_2658; // @[LZD.scala 39:25]
  wire [1:0] _T_2659; // @[Cat.scala 29:58]
  wire  _T_2660; // @[Shift.scala 12:21]
  wire  _T_2661; // @[Shift.scala 12:21]
  wire  _T_2662; // @[LZD.scala 49:16]
  wire  _T_2663; // @[LZD.scala 49:27]
  wire  _T_2664; // @[LZD.scala 49:25]
  wire  _T_2665; // @[LZD.scala 49:47]
  wire  _T_2666; // @[LZD.scala 49:59]
  wire  _T_2667; // @[LZD.scala 49:35]
  wire [2:0] _T_2669; // @[Cat.scala 29:58]
  wire [3:0] _T_2670; // @[LZD.scala 44:32]
  wire [1:0] _T_2671; // @[LZD.scala 43:32]
  wire  _T_2672; // @[LZD.scala 39:14]
  wire  _T_2673; // @[LZD.scala 39:21]
  wire  _T_2674; // @[LZD.scala 39:30]
  wire  _T_2675; // @[LZD.scala 39:27]
  wire  _T_2676; // @[LZD.scala 39:25]
  wire [1:0] _T_2677; // @[Cat.scala 29:58]
  wire [1:0] _T_2678; // @[LZD.scala 44:32]
  wire  _T_2679; // @[LZD.scala 39:14]
  wire  _T_2680; // @[LZD.scala 39:21]
  wire  _T_2681; // @[LZD.scala 39:30]
  wire  _T_2682; // @[LZD.scala 39:27]
  wire  _T_2683; // @[LZD.scala 39:25]
  wire [1:0] _T_2684; // @[Cat.scala 29:58]
  wire  _T_2685; // @[Shift.scala 12:21]
  wire  _T_2686; // @[Shift.scala 12:21]
  wire  _T_2687; // @[LZD.scala 49:16]
  wire  _T_2688; // @[LZD.scala 49:27]
  wire  _T_2689; // @[LZD.scala 49:25]
  wire  _T_2690; // @[LZD.scala 49:47]
  wire  _T_2691; // @[LZD.scala 49:59]
  wire  _T_2692; // @[LZD.scala 49:35]
  wire [2:0] _T_2694; // @[Cat.scala 29:58]
  wire  _T_2695; // @[Shift.scala 12:21]
  wire  _T_2696; // @[Shift.scala 12:21]
  wire  _T_2697; // @[LZD.scala 49:16]
  wire  _T_2698; // @[LZD.scala 49:27]
  wire  _T_2699; // @[LZD.scala 49:25]
  wire [1:0] _T_2700; // @[LZD.scala 49:47]
  wire [1:0] _T_2701; // @[LZD.scala 49:59]
  wire [1:0] _T_2702; // @[LZD.scala 49:35]
  wire [3:0] _T_2704; // @[Cat.scala 29:58]
  wire  _T_2705; // @[Shift.scala 12:21]
  wire  _T_2706; // @[Shift.scala 12:21]
  wire  _T_2707; // @[LZD.scala 49:16]
  wire  _T_2708; // @[LZD.scala 49:27]
  wire  _T_2709; // @[LZD.scala 49:25]
  wire [2:0] _T_2710; // @[LZD.scala 49:47]
  wire [2:0] _T_2711; // @[LZD.scala 49:59]
  wire [2:0] _T_2712; // @[LZD.scala 49:35]
  wire [4:0] _T_2714; // @[Cat.scala 29:58]
  wire [8:0] _T_2715; // @[LZD.scala 44:32]
  wire [7:0] _T_2716; // @[LZD.scala 43:32]
  wire [3:0] _T_2717; // @[LZD.scala 43:32]
  wire [1:0] _T_2718; // @[LZD.scala 43:32]
  wire  _T_2719; // @[LZD.scala 39:14]
  wire  _T_2720; // @[LZD.scala 39:21]
  wire  _T_2721; // @[LZD.scala 39:30]
  wire  _T_2722; // @[LZD.scala 39:27]
  wire  _T_2723; // @[LZD.scala 39:25]
  wire [1:0] _T_2724; // @[Cat.scala 29:58]
  wire [1:0] _T_2725; // @[LZD.scala 44:32]
  wire  _T_2726; // @[LZD.scala 39:14]
  wire  _T_2727; // @[LZD.scala 39:21]
  wire  _T_2728; // @[LZD.scala 39:30]
  wire  _T_2729; // @[LZD.scala 39:27]
  wire  _T_2730; // @[LZD.scala 39:25]
  wire [1:0] _T_2731; // @[Cat.scala 29:58]
  wire  _T_2732; // @[Shift.scala 12:21]
  wire  _T_2733; // @[Shift.scala 12:21]
  wire  _T_2734; // @[LZD.scala 49:16]
  wire  _T_2735; // @[LZD.scala 49:27]
  wire  _T_2736; // @[LZD.scala 49:25]
  wire  _T_2737; // @[LZD.scala 49:47]
  wire  _T_2738; // @[LZD.scala 49:59]
  wire  _T_2739; // @[LZD.scala 49:35]
  wire [2:0] _T_2741; // @[Cat.scala 29:58]
  wire [3:0] _T_2742; // @[LZD.scala 44:32]
  wire [1:0] _T_2743; // @[LZD.scala 43:32]
  wire  _T_2744; // @[LZD.scala 39:14]
  wire  _T_2745; // @[LZD.scala 39:21]
  wire  _T_2746; // @[LZD.scala 39:30]
  wire  _T_2747; // @[LZD.scala 39:27]
  wire  _T_2748; // @[LZD.scala 39:25]
  wire [1:0] _T_2749; // @[Cat.scala 29:58]
  wire [1:0] _T_2750; // @[LZD.scala 44:32]
  wire  _T_2751; // @[LZD.scala 39:14]
  wire  _T_2752; // @[LZD.scala 39:21]
  wire  _T_2753; // @[LZD.scala 39:30]
  wire  _T_2754; // @[LZD.scala 39:27]
  wire  _T_2755; // @[LZD.scala 39:25]
  wire [1:0] _T_2756; // @[Cat.scala 29:58]
  wire  _T_2757; // @[Shift.scala 12:21]
  wire  _T_2758; // @[Shift.scala 12:21]
  wire  _T_2759; // @[LZD.scala 49:16]
  wire  _T_2760; // @[LZD.scala 49:27]
  wire  _T_2761; // @[LZD.scala 49:25]
  wire  _T_2762; // @[LZD.scala 49:47]
  wire  _T_2763; // @[LZD.scala 49:59]
  wire  _T_2764; // @[LZD.scala 49:35]
  wire [2:0] _T_2766; // @[Cat.scala 29:58]
  wire  _T_2767; // @[Shift.scala 12:21]
  wire  _T_2768; // @[Shift.scala 12:21]
  wire  _T_2769; // @[LZD.scala 49:16]
  wire  _T_2770; // @[LZD.scala 49:27]
  wire  _T_2771; // @[LZD.scala 49:25]
  wire [1:0] _T_2772; // @[LZD.scala 49:47]
  wire [1:0] _T_2773; // @[LZD.scala 49:59]
  wire [1:0] _T_2774; // @[LZD.scala 49:35]
  wire [3:0] _T_2776; // @[Cat.scala 29:58]
  wire  _T_2777; // @[LZD.scala 44:32]
  wire  _T_2779; // @[Shift.scala 12:21]
  wire [2:0] _T_2782; // @[Cat.scala 29:58]
  wire [2:0] _T_2783; // @[LZD.scala 55:32]
  wire [2:0] _T_2784; // @[LZD.scala 55:20]
  wire [3:0] _T_2785; // @[Cat.scala 29:58]
  wire  _T_2786; // @[Shift.scala 12:21]
  wire [3:0] _T_2788; // @[LZD.scala 55:32]
  wire [3:0] _T_2789; // @[LZD.scala 55:20]
  wire [4:0] _T_2790; // @[Cat.scala 29:58]
  wire  _T_2791; // @[Shift.scala 12:21]
  wire [4:0] _T_2793; // @[LZD.scala 55:32]
  wire [4:0] _T_2794; // @[LZD.scala 55:20]
  wire  _T_2796; // @[Shift.scala 12:21]
  wire [7:0] _T_2799; // @[Cat.scala 29:58]
  wire [7:0] _T_2800; // @[LZD.scala 55:32]
  wire [7:0] _T_2801; // @[LZD.scala 55:20]
  wire [9:0] scaleBias; // @[Cat.scala 29:58]
  wire [9:0] _T_2802; // @[QuireToPosit.scala 61:53]
  wire [9:0] _T_2804; // @[QuireToPosit.scala 61:41]
  wire [9:0] realScale; // @[QuireToPosit.scala 61:41]
  wire  underflow; // @[QuireToPosit.scala 62:41]
  wire  overflow; // @[QuireToPosit.scala 63:35]
  wire [9:0] _T_2805; // @[Mux.scala 87:16]
  wire [9:0] _T_2806; // @[Mux.scala 87:16]
  wire  _T_2807; // @[Abs.scala 10:21]
  wire [9:0] _T_2809; // @[Bitwise.scala 71:12]
  wire [9:0] _T_2810; // @[Abs.scala 10:31]
  wire [9:0] _T_2811; // @[Abs.scala 10:26]
  wire [9:0] _GEN_2; // @[Abs.scala 10:39]
  wire [9:0] absRealScale; // @[Abs.scala 10:39]
  wire  _T_2814; // @[Shift.scala 16:24]
  wire [8:0] _T_2815; // @[Shift.scala 17:37]
  wire  _T_2816; // @[Shift.scala 12:21]
  wire [57:0] _T_2817; // @[Shift.scala 64:52]
  wire [313:0] _T_2819; // @[Cat.scala 29:58]
  wire [313:0] _T_2820; // @[Shift.scala 64:27]
  wire [7:0] _T_2821; // @[Shift.scala 66:70]
  wire  _T_2822; // @[Shift.scala 12:21]
  wire [185:0] _T_2823; // @[Shift.scala 64:52]
  wire [313:0] _T_2825; // @[Cat.scala 29:58]
  wire [313:0] _T_2826; // @[Shift.scala 64:27]
  wire [6:0] _T_2827; // @[Shift.scala 66:70]
  wire  _T_2828; // @[Shift.scala 12:21]
  wire [249:0] _T_2829; // @[Shift.scala 64:52]
  wire [313:0] _T_2831; // @[Cat.scala 29:58]
  wire [313:0] _T_2832; // @[Shift.scala 64:27]
  wire [5:0] _T_2833; // @[Shift.scala 66:70]
  wire  _T_2834; // @[Shift.scala 12:21]
  wire [281:0] _T_2835; // @[Shift.scala 64:52]
  wire [313:0] _T_2837; // @[Cat.scala 29:58]
  wire [313:0] _T_2838; // @[Shift.scala 64:27]
  wire [4:0] _T_2839; // @[Shift.scala 66:70]
  wire  _T_2840; // @[Shift.scala 12:21]
  wire [297:0] _T_2841; // @[Shift.scala 64:52]
  wire [313:0] _T_2843; // @[Cat.scala 29:58]
  wire [313:0] _T_2844; // @[Shift.scala 64:27]
  wire [3:0] _T_2845; // @[Shift.scala 66:70]
  wire  _T_2846; // @[Shift.scala 12:21]
  wire [305:0] _T_2847; // @[Shift.scala 64:52]
  wire [313:0] _T_2849; // @[Cat.scala 29:58]
  wire [313:0] _T_2850; // @[Shift.scala 64:27]
  wire [2:0] _T_2851; // @[Shift.scala 66:70]
  wire  _T_2852; // @[Shift.scala 12:21]
  wire [309:0] _T_2853; // @[Shift.scala 64:52]
  wire [313:0] _T_2855; // @[Cat.scala 29:58]
  wire [313:0] _T_2856; // @[Shift.scala 64:27]
  wire [1:0] _T_2857; // @[Shift.scala 66:70]
  wire  _T_2858; // @[Shift.scala 12:21]
  wire [311:0] _T_2859; // @[Shift.scala 64:52]
  wire [313:0] _T_2861; // @[Cat.scala 29:58]
  wire [313:0] _T_2862; // @[Shift.scala 64:27]
  wire  _T_2863; // @[Shift.scala 66:70]
  wire [312:0] _T_2865; // @[Shift.scala 64:52]
  wire [313:0] _T_2866; // @[Cat.scala 29:58]
  wire [313:0] _T_2867; // @[Shift.scala 64:27]
  wire [313:0] quireLeftShift; // @[Shift.scala 16:10]
  wire [57:0] _T_2872; // @[Shift.scala 77:66]
  wire [313:0] _T_2873; // @[Cat.scala 29:58]
  wire [313:0] _T_2874; // @[Shift.scala 77:22]
  wire [185:0] _T_2878; // @[Shift.scala 77:66]
  wire [313:0] _T_2879; // @[Cat.scala 29:58]
  wire [313:0] _T_2880; // @[Shift.scala 77:22]
  wire [249:0] _T_2884; // @[Shift.scala 77:66]
  wire [313:0] _T_2885; // @[Cat.scala 29:58]
  wire [313:0] _T_2886; // @[Shift.scala 77:22]
  wire [281:0] _T_2890; // @[Shift.scala 77:66]
  wire [313:0] _T_2891; // @[Cat.scala 29:58]
  wire [313:0] _T_2892; // @[Shift.scala 77:22]
  wire [297:0] _T_2896; // @[Shift.scala 77:66]
  wire [313:0] _T_2897; // @[Cat.scala 29:58]
  wire [313:0] _T_2898; // @[Shift.scala 77:22]
  wire [305:0] _T_2902; // @[Shift.scala 77:66]
  wire [313:0] _T_2903; // @[Cat.scala 29:58]
  wire [313:0] _T_2904; // @[Shift.scala 77:22]
  wire [309:0] _T_2908; // @[Shift.scala 77:66]
  wire [313:0] _T_2909; // @[Cat.scala 29:58]
  wire [313:0] _T_2910; // @[Shift.scala 77:22]
  wire [311:0] _T_2914; // @[Shift.scala 77:66]
  wire [313:0] _T_2915; // @[Cat.scala 29:58]
  wire [313:0] _T_2916; // @[Shift.scala 77:22]
  wire [312:0] _T_2919; // @[Shift.scala 77:66]
  wire [313:0] _T_2920; // @[Cat.scala 29:58]
  wire [313:0] _T_2921; // @[Shift.scala 77:22]
  wire [313:0] quireRightShift; // @[Shift.scala 27:10]
  wire [14:0] _T_2923; // @[QuireToPosit.scala 89:49]
  wire [12:0] _T_2924; // @[QuireToPosit.scala 90:127]
  wire  _T_2925; // @[QuireToPosit.scala 90:154]
  wire [15:0] realFGRSTmp1; // @[Cat.scala 29:58]
  wire [14:0] _T_2926; // @[QuireToPosit.scala 91:50]
  wire [12:0] _T_2927; // @[QuireToPosit.scala 92:128]
  wire  _T_2928; // @[QuireToPosit.scala 92:155]
  wire [15:0] realFGRSTmp2; // @[Cat.scala 29:58]
  wire [15:0] realFGRS; // @[QuireToPosit.scala 93:34]
  wire [12:0] outRawFloat_fraction; // @[QuireToPosit.scala 95:46]
  wire [2:0] outRawFloat_grs; // @[QuireToPosit.scala 96:46]
  wire [4:0] _GEN_3; // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  wire [4:0] outRawFloat_scale; // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  wire  _T_2934; // @[convert.scala 49:36]
  wire [4:0] _T_2936; // @[convert.scala 50:36]
  wire [4:0] _T_2937; // @[convert.scala 50:36]
  wire [4:0] _T_2938; // @[convert.scala 50:28]
  wire  _T_2939; // @[convert.scala 51:31]
  wire  _T_2940; // @[convert.scala 53:34]
  wire [17:0] _T_2943; // @[Cat.scala 29:58]
  wire [4:0] _T_2944; // @[Shift.scala 39:17]
  wire  _T_2945; // @[Shift.scala 39:24]
  wire [1:0] _T_2947; // @[Shift.scala 90:30]
  wire [15:0] _T_2948; // @[Shift.scala 90:48]
  wire  _T_2949; // @[Shift.scala 90:57]
  wire [1:0] _GEN_4; // @[Shift.scala 90:39]
  wire [1:0] _T_2950; // @[Shift.scala 90:39]
  wire  _T_2951; // @[Shift.scala 12:21]
  wire  _T_2952; // @[Shift.scala 12:21]
  wire [15:0] _T_2954; // @[Bitwise.scala 71:12]
  wire [17:0] _T_2955; // @[Cat.scala 29:58]
  wire [17:0] _T_2956; // @[Shift.scala 91:22]
  wire [3:0] _T_2957; // @[Shift.scala 92:77]
  wire [9:0] _T_2958; // @[Shift.scala 90:30]
  wire [7:0] _T_2959; // @[Shift.scala 90:48]
  wire  _T_2960; // @[Shift.scala 90:57]
  wire [9:0] _GEN_5; // @[Shift.scala 90:39]
  wire [9:0] _T_2961; // @[Shift.scala 90:39]
  wire  _T_2962; // @[Shift.scala 12:21]
  wire  _T_2963; // @[Shift.scala 12:21]
  wire [7:0] _T_2965; // @[Bitwise.scala 71:12]
  wire [17:0] _T_2966; // @[Cat.scala 29:58]
  wire [17:0] _T_2967; // @[Shift.scala 91:22]
  wire [2:0] _T_2968; // @[Shift.scala 92:77]
  wire [13:0] _T_2969; // @[Shift.scala 90:30]
  wire [3:0] _T_2970; // @[Shift.scala 90:48]
  wire  _T_2971; // @[Shift.scala 90:57]
  wire [13:0] _GEN_6; // @[Shift.scala 90:39]
  wire [13:0] _T_2972; // @[Shift.scala 90:39]
  wire  _T_2973; // @[Shift.scala 12:21]
  wire  _T_2974; // @[Shift.scala 12:21]
  wire [3:0] _T_2976; // @[Bitwise.scala 71:12]
  wire [17:0] _T_2977; // @[Cat.scala 29:58]
  wire [17:0] _T_2978; // @[Shift.scala 91:22]
  wire [1:0] _T_2979; // @[Shift.scala 92:77]
  wire [15:0] _T_2980; // @[Shift.scala 90:30]
  wire [1:0] _T_2981; // @[Shift.scala 90:48]
  wire  _T_2982; // @[Shift.scala 90:57]
  wire [15:0] _GEN_7; // @[Shift.scala 90:39]
  wire [15:0] _T_2983; // @[Shift.scala 90:39]
  wire  _T_2984; // @[Shift.scala 12:21]
  wire  _T_2985; // @[Shift.scala 12:21]
  wire [1:0] _T_2987; // @[Bitwise.scala 71:12]
  wire [17:0] _T_2988; // @[Cat.scala 29:58]
  wire [17:0] _T_2989; // @[Shift.scala 91:22]
  wire  _T_2990; // @[Shift.scala 92:77]
  wire [16:0] _T_2991; // @[Shift.scala 90:30]
  wire  _T_2992; // @[Shift.scala 90:48]
  wire [16:0] _GEN_8; // @[Shift.scala 90:39]
  wire [16:0] _T_2994; // @[Shift.scala 90:39]
  wire  _T_2996; // @[Shift.scala 12:21]
  wire [17:0] _T_2997; // @[Cat.scala 29:58]
  wire [17:0] _T_2998; // @[Shift.scala 91:22]
  wire [17:0] _T_3001; // @[Bitwise.scala 71:12]
  wire [17:0] _T_3002; // @[Shift.scala 39:10]
  wire  _T_3003; // @[convert.scala 55:31]
  wire  _T_3004; // @[convert.scala 56:31]
  wire  _T_3005; // @[convert.scala 57:31]
  wire  _T_3006; // @[convert.scala 58:31]
  wire [14:0] _T_3007; // @[convert.scala 59:69]
  wire  _T_3008; // @[convert.scala 59:81]
  wire  _T_3009; // @[convert.scala 59:50]
  wire  _T_3011; // @[convert.scala 60:81]
  wire  _T_3012; // @[convert.scala 61:44]
  wire  _T_3013; // @[convert.scala 61:52]
  wire  _T_3014; // @[convert.scala 61:36]
  wire  _T_3015; // @[convert.scala 62:63]
  wire  _T_3016; // @[convert.scala 62:103]
  wire  _T_3017; // @[convert.scala 62:60]
  wire [14:0] _GEN_9; // @[convert.scala 63:56]
  wire [14:0] _T_3020; // @[convert.scala 63:56]
  wire [15:0] _T_3021; // @[Cat.scala 29:58]
  reg  _T_3025; // @[Valid.scala 117:22]
  reg [31:0] _RAND_0;
  reg [15:0] _T_3029; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  assign _T = io_quireIn[312:0]; // @[QuireToPosit.scala 47:43]
  assign _T_1 = _T != 313'h0; // @[QuireToPosit.scala 47:47]
  assign tailIsZero = ~ _T_1; // @[QuireToPosit.scala 47:27]
  assign _T_2 = io_quireIn[313:313]; // @[QuireToPosit.scala 49:45]
  assign outRawFloat_isNaR = _T_2 & tailIsZero; // @[QuireToPosit.scala 49:49]
  assign _T_5 = ~ _T_2; // @[QuireToPosit.scala 50:31]
  assign outRawFloat_isZero = _T_5 & tailIsZero; // @[QuireToPosit.scala 50:51]
  assign _T_8 = io_quireIn[313:1]; // @[QuireToPosit.scala 58:41]
  assign _T_9 = io_quireIn[312:0]; // @[QuireToPosit.scala 58:68]
  assign quireXOR = _T_8 ^ _T_9; // @[QuireToPosit.scala 58:56]
  assign _T_10 = quireXOR[312:57]; // @[LZD.scala 43:32]
  assign _T_11 = _T_10[255:128]; // @[LZD.scala 43:32]
  assign _T_12 = _T_11[127:64]; // @[LZD.scala 43:32]
  assign _T_13 = _T_12[63:32]; // @[LZD.scala 43:32]
  assign _T_14 = _T_13[31:16]; // @[LZD.scala 43:32]
  assign _T_15 = _T_14[15:8]; // @[LZD.scala 43:32]
  assign _T_16 = _T_15[7:4]; // @[LZD.scala 43:32]
  assign _T_17 = _T_16[3:2]; // @[LZD.scala 43:32]
  assign _T_18 = _T_17 != 2'h0; // @[LZD.scala 39:14]
  assign _T_19 = _T_17[1]; // @[LZD.scala 39:21]
  assign _T_20 = _T_17[0]; // @[LZD.scala 39:30]
  assign _T_21 = ~ _T_20; // @[LZD.scala 39:27]
  assign _T_22 = _T_19 | _T_21; // @[LZD.scala 39:25]
  assign _T_23 = {_T_18,_T_22}; // @[Cat.scala 29:58]
  assign _T_24 = _T_16[1:0]; // @[LZD.scala 44:32]
  assign _T_25 = _T_24 != 2'h0; // @[LZD.scala 39:14]
  assign _T_26 = _T_24[1]; // @[LZD.scala 39:21]
  assign _T_27 = _T_24[0]; // @[LZD.scala 39:30]
  assign _T_28 = ~ _T_27; // @[LZD.scala 39:27]
  assign _T_29 = _T_26 | _T_28; // @[LZD.scala 39:25]
  assign _T_30 = {_T_25,_T_29}; // @[Cat.scala 29:58]
  assign _T_31 = _T_23[1]; // @[Shift.scala 12:21]
  assign _T_32 = _T_30[1]; // @[Shift.scala 12:21]
  assign _T_33 = _T_31 | _T_32; // @[LZD.scala 49:16]
  assign _T_34 = ~ _T_32; // @[LZD.scala 49:27]
  assign _T_35 = _T_31 | _T_34; // @[LZD.scala 49:25]
  assign _T_36 = _T_23[0:0]; // @[LZD.scala 49:47]
  assign _T_37 = _T_30[0:0]; // @[LZD.scala 49:59]
  assign _T_38 = _T_31 ? _T_36 : _T_37; // @[LZD.scala 49:35]
  assign _T_40 = {_T_33,_T_35,_T_38}; // @[Cat.scala 29:58]
  assign _T_41 = _T_15[3:0]; // @[LZD.scala 44:32]
  assign _T_42 = _T_41[3:2]; // @[LZD.scala 43:32]
  assign _T_43 = _T_42 != 2'h0; // @[LZD.scala 39:14]
  assign _T_44 = _T_42[1]; // @[LZD.scala 39:21]
  assign _T_45 = _T_42[0]; // @[LZD.scala 39:30]
  assign _T_46 = ~ _T_45; // @[LZD.scala 39:27]
  assign _T_47 = _T_44 | _T_46; // @[LZD.scala 39:25]
  assign _T_48 = {_T_43,_T_47}; // @[Cat.scala 29:58]
  assign _T_49 = _T_41[1:0]; // @[LZD.scala 44:32]
  assign _T_50 = _T_49 != 2'h0; // @[LZD.scala 39:14]
  assign _T_51 = _T_49[1]; // @[LZD.scala 39:21]
  assign _T_52 = _T_49[0]; // @[LZD.scala 39:30]
  assign _T_53 = ~ _T_52; // @[LZD.scala 39:27]
  assign _T_54 = _T_51 | _T_53; // @[LZD.scala 39:25]
  assign _T_55 = {_T_50,_T_54}; // @[Cat.scala 29:58]
  assign _T_56 = _T_48[1]; // @[Shift.scala 12:21]
  assign _T_57 = _T_55[1]; // @[Shift.scala 12:21]
  assign _T_58 = _T_56 | _T_57; // @[LZD.scala 49:16]
  assign _T_59 = ~ _T_57; // @[LZD.scala 49:27]
  assign _T_60 = _T_56 | _T_59; // @[LZD.scala 49:25]
  assign _T_61 = _T_48[0:0]; // @[LZD.scala 49:47]
  assign _T_62 = _T_55[0:0]; // @[LZD.scala 49:59]
  assign _T_63 = _T_56 ? _T_61 : _T_62; // @[LZD.scala 49:35]
  assign _T_65 = {_T_58,_T_60,_T_63}; // @[Cat.scala 29:58]
  assign _T_66 = _T_40[2]; // @[Shift.scala 12:21]
  assign _T_67 = _T_65[2]; // @[Shift.scala 12:21]
  assign _T_68 = _T_66 | _T_67; // @[LZD.scala 49:16]
  assign _T_69 = ~ _T_67; // @[LZD.scala 49:27]
  assign _T_70 = _T_66 | _T_69; // @[LZD.scala 49:25]
  assign _T_71 = _T_40[1:0]; // @[LZD.scala 49:47]
  assign _T_72 = _T_65[1:0]; // @[LZD.scala 49:59]
  assign _T_73 = _T_66 ? _T_71 : _T_72; // @[LZD.scala 49:35]
  assign _T_75 = {_T_68,_T_70,_T_73}; // @[Cat.scala 29:58]
  assign _T_76 = _T_14[7:0]; // @[LZD.scala 44:32]
  assign _T_77 = _T_76[7:4]; // @[LZD.scala 43:32]
  assign _T_78 = _T_77[3:2]; // @[LZD.scala 43:32]
  assign _T_79 = _T_78 != 2'h0; // @[LZD.scala 39:14]
  assign _T_80 = _T_78[1]; // @[LZD.scala 39:21]
  assign _T_81 = _T_78[0]; // @[LZD.scala 39:30]
  assign _T_82 = ~ _T_81; // @[LZD.scala 39:27]
  assign _T_83 = _T_80 | _T_82; // @[LZD.scala 39:25]
  assign _T_84 = {_T_79,_T_83}; // @[Cat.scala 29:58]
  assign _T_85 = _T_77[1:0]; // @[LZD.scala 44:32]
  assign _T_86 = _T_85 != 2'h0; // @[LZD.scala 39:14]
  assign _T_87 = _T_85[1]; // @[LZD.scala 39:21]
  assign _T_88 = _T_85[0]; // @[LZD.scala 39:30]
  assign _T_89 = ~ _T_88; // @[LZD.scala 39:27]
  assign _T_90 = _T_87 | _T_89; // @[LZD.scala 39:25]
  assign _T_91 = {_T_86,_T_90}; // @[Cat.scala 29:58]
  assign _T_92 = _T_84[1]; // @[Shift.scala 12:21]
  assign _T_93 = _T_91[1]; // @[Shift.scala 12:21]
  assign _T_94 = _T_92 | _T_93; // @[LZD.scala 49:16]
  assign _T_95 = ~ _T_93; // @[LZD.scala 49:27]
  assign _T_96 = _T_92 | _T_95; // @[LZD.scala 49:25]
  assign _T_97 = _T_84[0:0]; // @[LZD.scala 49:47]
  assign _T_98 = _T_91[0:0]; // @[LZD.scala 49:59]
  assign _T_99 = _T_92 ? _T_97 : _T_98; // @[LZD.scala 49:35]
  assign _T_101 = {_T_94,_T_96,_T_99}; // @[Cat.scala 29:58]
  assign _T_102 = _T_76[3:0]; // @[LZD.scala 44:32]
  assign _T_103 = _T_102[3:2]; // @[LZD.scala 43:32]
  assign _T_104 = _T_103 != 2'h0; // @[LZD.scala 39:14]
  assign _T_105 = _T_103[1]; // @[LZD.scala 39:21]
  assign _T_106 = _T_103[0]; // @[LZD.scala 39:30]
  assign _T_107 = ~ _T_106; // @[LZD.scala 39:27]
  assign _T_108 = _T_105 | _T_107; // @[LZD.scala 39:25]
  assign _T_109 = {_T_104,_T_108}; // @[Cat.scala 29:58]
  assign _T_110 = _T_102[1:0]; // @[LZD.scala 44:32]
  assign _T_111 = _T_110 != 2'h0; // @[LZD.scala 39:14]
  assign _T_112 = _T_110[1]; // @[LZD.scala 39:21]
  assign _T_113 = _T_110[0]; // @[LZD.scala 39:30]
  assign _T_114 = ~ _T_113; // @[LZD.scala 39:27]
  assign _T_115 = _T_112 | _T_114; // @[LZD.scala 39:25]
  assign _T_116 = {_T_111,_T_115}; // @[Cat.scala 29:58]
  assign _T_117 = _T_109[1]; // @[Shift.scala 12:21]
  assign _T_118 = _T_116[1]; // @[Shift.scala 12:21]
  assign _T_119 = _T_117 | _T_118; // @[LZD.scala 49:16]
  assign _T_120 = ~ _T_118; // @[LZD.scala 49:27]
  assign _T_121 = _T_117 | _T_120; // @[LZD.scala 49:25]
  assign _T_122 = _T_109[0:0]; // @[LZD.scala 49:47]
  assign _T_123 = _T_116[0:0]; // @[LZD.scala 49:59]
  assign _T_124 = _T_117 ? _T_122 : _T_123; // @[LZD.scala 49:35]
  assign _T_126 = {_T_119,_T_121,_T_124}; // @[Cat.scala 29:58]
  assign _T_127 = _T_101[2]; // @[Shift.scala 12:21]
  assign _T_128 = _T_126[2]; // @[Shift.scala 12:21]
  assign _T_129 = _T_127 | _T_128; // @[LZD.scala 49:16]
  assign _T_130 = ~ _T_128; // @[LZD.scala 49:27]
  assign _T_131 = _T_127 | _T_130; // @[LZD.scala 49:25]
  assign _T_132 = _T_101[1:0]; // @[LZD.scala 49:47]
  assign _T_133 = _T_126[1:0]; // @[LZD.scala 49:59]
  assign _T_134 = _T_127 ? _T_132 : _T_133; // @[LZD.scala 49:35]
  assign _T_136 = {_T_129,_T_131,_T_134}; // @[Cat.scala 29:58]
  assign _T_137 = _T_75[3]; // @[Shift.scala 12:21]
  assign _T_138 = _T_136[3]; // @[Shift.scala 12:21]
  assign _T_139 = _T_137 | _T_138; // @[LZD.scala 49:16]
  assign _T_140 = ~ _T_138; // @[LZD.scala 49:27]
  assign _T_141 = _T_137 | _T_140; // @[LZD.scala 49:25]
  assign _T_142 = _T_75[2:0]; // @[LZD.scala 49:47]
  assign _T_143 = _T_136[2:0]; // @[LZD.scala 49:59]
  assign _T_144 = _T_137 ? _T_142 : _T_143; // @[LZD.scala 49:35]
  assign _T_146 = {_T_139,_T_141,_T_144}; // @[Cat.scala 29:58]
  assign _T_147 = _T_13[15:0]; // @[LZD.scala 44:32]
  assign _T_148 = _T_147[15:8]; // @[LZD.scala 43:32]
  assign _T_149 = _T_148[7:4]; // @[LZD.scala 43:32]
  assign _T_150 = _T_149[3:2]; // @[LZD.scala 43:32]
  assign _T_151 = _T_150 != 2'h0; // @[LZD.scala 39:14]
  assign _T_152 = _T_150[1]; // @[LZD.scala 39:21]
  assign _T_153 = _T_150[0]; // @[LZD.scala 39:30]
  assign _T_154 = ~ _T_153; // @[LZD.scala 39:27]
  assign _T_155 = _T_152 | _T_154; // @[LZD.scala 39:25]
  assign _T_156 = {_T_151,_T_155}; // @[Cat.scala 29:58]
  assign _T_157 = _T_149[1:0]; // @[LZD.scala 44:32]
  assign _T_158 = _T_157 != 2'h0; // @[LZD.scala 39:14]
  assign _T_159 = _T_157[1]; // @[LZD.scala 39:21]
  assign _T_160 = _T_157[0]; // @[LZD.scala 39:30]
  assign _T_161 = ~ _T_160; // @[LZD.scala 39:27]
  assign _T_162 = _T_159 | _T_161; // @[LZD.scala 39:25]
  assign _T_163 = {_T_158,_T_162}; // @[Cat.scala 29:58]
  assign _T_164 = _T_156[1]; // @[Shift.scala 12:21]
  assign _T_165 = _T_163[1]; // @[Shift.scala 12:21]
  assign _T_166 = _T_164 | _T_165; // @[LZD.scala 49:16]
  assign _T_167 = ~ _T_165; // @[LZD.scala 49:27]
  assign _T_168 = _T_164 | _T_167; // @[LZD.scala 49:25]
  assign _T_169 = _T_156[0:0]; // @[LZD.scala 49:47]
  assign _T_170 = _T_163[0:0]; // @[LZD.scala 49:59]
  assign _T_171 = _T_164 ? _T_169 : _T_170; // @[LZD.scala 49:35]
  assign _T_173 = {_T_166,_T_168,_T_171}; // @[Cat.scala 29:58]
  assign _T_174 = _T_148[3:0]; // @[LZD.scala 44:32]
  assign _T_175 = _T_174[3:2]; // @[LZD.scala 43:32]
  assign _T_176 = _T_175 != 2'h0; // @[LZD.scala 39:14]
  assign _T_177 = _T_175[1]; // @[LZD.scala 39:21]
  assign _T_178 = _T_175[0]; // @[LZD.scala 39:30]
  assign _T_179 = ~ _T_178; // @[LZD.scala 39:27]
  assign _T_180 = _T_177 | _T_179; // @[LZD.scala 39:25]
  assign _T_181 = {_T_176,_T_180}; // @[Cat.scala 29:58]
  assign _T_182 = _T_174[1:0]; // @[LZD.scala 44:32]
  assign _T_183 = _T_182 != 2'h0; // @[LZD.scala 39:14]
  assign _T_184 = _T_182[1]; // @[LZD.scala 39:21]
  assign _T_185 = _T_182[0]; // @[LZD.scala 39:30]
  assign _T_186 = ~ _T_185; // @[LZD.scala 39:27]
  assign _T_187 = _T_184 | _T_186; // @[LZD.scala 39:25]
  assign _T_188 = {_T_183,_T_187}; // @[Cat.scala 29:58]
  assign _T_189 = _T_181[1]; // @[Shift.scala 12:21]
  assign _T_190 = _T_188[1]; // @[Shift.scala 12:21]
  assign _T_191 = _T_189 | _T_190; // @[LZD.scala 49:16]
  assign _T_192 = ~ _T_190; // @[LZD.scala 49:27]
  assign _T_193 = _T_189 | _T_192; // @[LZD.scala 49:25]
  assign _T_194 = _T_181[0:0]; // @[LZD.scala 49:47]
  assign _T_195 = _T_188[0:0]; // @[LZD.scala 49:59]
  assign _T_196 = _T_189 ? _T_194 : _T_195; // @[LZD.scala 49:35]
  assign _T_198 = {_T_191,_T_193,_T_196}; // @[Cat.scala 29:58]
  assign _T_199 = _T_173[2]; // @[Shift.scala 12:21]
  assign _T_200 = _T_198[2]; // @[Shift.scala 12:21]
  assign _T_201 = _T_199 | _T_200; // @[LZD.scala 49:16]
  assign _T_202 = ~ _T_200; // @[LZD.scala 49:27]
  assign _T_203 = _T_199 | _T_202; // @[LZD.scala 49:25]
  assign _T_204 = _T_173[1:0]; // @[LZD.scala 49:47]
  assign _T_205 = _T_198[1:0]; // @[LZD.scala 49:59]
  assign _T_206 = _T_199 ? _T_204 : _T_205; // @[LZD.scala 49:35]
  assign _T_208 = {_T_201,_T_203,_T_206}; // @[Cat.scala 29:58]
  assign _T_209 = _T_147[7:0]; // @[LZD.scala 44:32]
  assign _T_210 = _T_209[7:4]; // @[LZD.scala 43:32]
  assign _T_211 = _T_210[3:2]; // @[LZD.scala 43:32]
  assign _T_212 = _T_211 != 2'h0; // @[LZD.scala 39:14]
  assign _T_213 = _T_211[1]; // @[LZD.scala 39:21]
  assign _T_214 = _T_211[0]; // @[LZD.scala 39:30]
  assign _T_215 = ~ _T_214; // @[LZD.scala 39:27]
  assign _T_216 = _T_213 | _T_215; // @[LZD.scala 39:25]
  assign _T_217 = {_T_212,_T_216}; // @[Cat.scala 29:58]
  assign _T_218 = _T_210[1:0]; // @[LZD.scala 44:32]
  assign _T_219 = _T_218 != 2'h0; // @[LZD.scala 39:14]
  assign _T_220 = _T_218[1]; // @[LZD.scala 39:21]
  assign _T_221 = _T_218[0]; // @[LZD.scala 39:30]
  assign _T_222 = ~ _T_221; // @[LZD.scala 39:27]
  assign _T_223 = _T_220 | _T_222; // @[LZD.scala 39:25]
  assign _T_224 = {_T_219,_T_223}; // @[Cat.scala 29:58]
  assign _T_225 = _T_217[1]; // @[Shift.scala 12:21]
  assign _T_226 = _T_224[1]; // @[Shift.scala 12:21]
  assign _T_227 = _T_225 | _T_226; // @[LZD.scala 49:16]
  assign _T_228 = ~ _T_226; // @[LZD.scala 49:27]
  assign _T_229 = _T_225 | _T_228; // @[LZD.scala 49:25]
  assign _T_230 = _T_217[0:0]; // @[LZD.scala 49:47]
  assign _T_231 = _T_224[0:0]; // @[LZD.scala 49:59]
  assign _T_232 = _T_225 ? _T_230 : _T_231; // @[LZD.scala 49:35]
  assign _T_234 = {_T_227,_T_229,_T_232}; // @[Cat.scala 29:58]
  assign _T_235 = _T_209[3:0]; // @[LZD.scala 44:32]
  assign _T_236 = _T_235[3:2]; // @[LZD.scala 43:32]
  assign _T_237 = _T_236 != 2'h0; // @[LZD.scala 39:14]
  assign _T_238 = _T_236[1]; // @[LZD.scala 39:21]
  assign _T_239 = _T_236[0]; // @[LZD.scala 39:30]
  assign _T_240 = ~ _T_239; // @[LZD.scala 39:27]
  assign _T_241 = _T_238 | _T_240; // @[LZD.scala 39:25]
  assign _T_242 = {_T_237,_T_241}; // @[Cat.scala 29:58]
  assign _T_243 = _T_235[1:0]; // @[LZD.scala 44:32]
  assign _T_244 = _T_243 != 2'h0; // @[LZD.scala 39:14]
  assign _T_245 = _T_243[1]; // @[LZD.scala 39:21]
  assign _T_246 = _T_243[0]; // @[LZD.scala 39:30]
  assign _T_247 = ~ _T_246; // @[LZD.scala 39:27]
  assign _T_248 = _T_245 | _T_247; // @[LZD.scala 39:25]
  assign _T_249 = {_T_244,_T_248}; // @[Cat.scala 29:58]
  assign _T_250 = _T_242[1]; // @[Shift.scala 12:21]
  assign _T_251 = _T_249[1]; // @[Shift.scala 12:21]
  assign _T_252 = _T_250 | _T_251; // @[LZD.scala 49:16]
  assign _T_253 = ~ _T_251; // @[LZD.scala 49:27]
  assign _T_254 = _T_250 | _T_253; // @[LZD.scala 49:25]
  assign _T_255 = _T_242[0:0]; // @[LZD.scala 49:47]
  assign _T_256 = _T_249[0:0]; // @[LZD.scala 49:59]
  assign _T_257 = _T_250 ? _T_255 : _T_256; // @[LZD.scala 49:35]
  assign _T_259 = {_T_252,_T_254,_T_257}; // @[Cat.scala 29:58]
  assign _T_260 = _T_234[2]; // @[Shift.scala 12:21]
  assign _T_261 = _T_259[2]; // @[Shift.scala 12:21]
  assign _T_262 = _T_260 | _T_261; // @[LZD.scala 49:16]
  assign _T_263 = ~ _T_261; // @[LZD.scala 49:27]
  assign _T_264 = _T_260 | _T_263; // @[LZD.scala 49:25]
  assign _T_265 = _T_234[1:0]; // @[LZD.scala 49:47]
  assign _T_266 = _T_259[1:0]; // @[LZD.scala 49:59]
  assign _T_267 = _T_260 ? _T_265 : _T_266; // @[LZD.scala 49:35]
  assign _T_269 = {_T_262,_T_264,_T_267}; // @[Cat.scala 29:58]
  assign _T_270 = _T_208[3]; // @[Shift.scala 12:21]
  assign _T_271 = _T_269[3]; // @[Shift.scala 12:21]
  assign _T_272 = _T_270 | _T_271; // @[LZD.scala 49:16]
  assign _T_273 = ~ _T_271; // @[LZD.scala 49:27]
  assign _T_274 = _T_270 | _T_273; // @[LZD.scala 49:25]
  assign _T_275 = _T_208[2:0]; // @[LZD.scala 49:47]
  assign _T_276 = _T_269[2:0]; // @[LZD.scala 49:59]
  assign _T_277 = _T_270 ? _T_275 : _T_276; // @[LZD.scala 49:35]
  assign _T_279 = {_T_272,_T_274,_T_277}; // @[Cat.scala 29:58]
  assign _T_280 = _T_146[4]; // @[Shift.scala 12:21]
  assign _T_281 = _T_279[4]; // @[Shift.scala 12:21]
  assign _T_282 = _T_280 | _T_281; // @[LZD.scala 49:16]
  assign _T_283 = ~ _T_281; // @[LZD.scala 49:27]
  assign _T_284 = _T_280 | _T_283; // @[LZD.scala 49:25]
  assign _T_285 = _T_146[3:0]; // @[LZD.scala 49:47]
  assign _T_286 = _T_279[3:0]; // @[LZD.scala 49:59]
  assign _T_287 = _T_280 ? _T_285 : _T_286; // @[LZD.scala 49:35]
  assign _T_289 = {_T_282,_T_284,_T_287}; // @[Cat.scala 29:58]
  assign _T_290 = _T_12[31:0]; // @[LZD.scala 44:32]
  assign _T_291 = _T_290[31:16]; // @[LZD.scala 43:32]
  assign _T_292 = _T_291[15:8]; // @[LZD.scala 43:32]
  assign _T_293 = _T_292[7:4]; // @[LZD.scala 43:32]
  assign _T_294 = _T_293[3:2]; // @[LZD.scala 43:32]
  assign _T_295 = _T_294 != 2'h0; // @[LZD.scala 39:14]
  assign _T_296 = _T_294[1]; // @[LZD.scala 39:21]
  assign _T_297 = _T_294[0]; // @[LZD.scala 39:30]
  assign _T_298 = ~ _T_297; // @[LZD.scala 39:27]
  assign _T_299 = _T_296 | _T_298; // @[LZD.scala 39:25]
  assign _T_300 = {_T_295,_T_299}; // @[Cat.scala 29:58]
  assign _T_301 = _T_293[1:0]; // @[LZD.scala 44:32]
  assign _T_302 = _T_301 != 2'h0; // @[LZD.scala 39:14]
  assign _T_303 = _T_301[1]; // @[LZD.scala 39:21]
  assign _T_304 = _T_301[0]; // @[LZD.scala 39:30]
  assign _T_305 = ~ _T_304; // @[LZD.scala 39:27]
  assign _T_306 = _T_303 | _T_305; // @[LZD.scala 39:25]
  assign _T_307 = {_T_302,_T_306}; // @[Cat.scala 29:58]
  assign _T_308 = _T_300[1]; // @[Shift.scala 12:21]
  assign _T_309 = _T_307[1]; // @[Shift.scala 12:21]
  assign _T_310 = _T_308 | _T_309; // @[LZD.scala 49:16]
  assign _T_311 = ~ _T_309; // @[LZD.scala 49:27]
  assign _T_312 = _T_308 | _T_311; // @[LZD.scala 49:25]
  assign _T_313 = _T_300[0:0]; // @[LZD.scala 49:47]
  assign _T_314 = _T_307[0:0]; // @[LZD.scala 49:59]
  assign _T_315 = _T_308 ? _T_313 : _T_314; // @[LZD.scala 49:35]
  assign _T_317 = {_T_310,_T_312,_T_315}; // @[Cat.scala 29:58]
  assign _T_318 = _T_292[3:0]; // @[LZD.scala 44:32]
  assign _T_319 = _T_318[3:2]; // @[LZD.scala 43:32]
  assign _T_320 = _T_319 != 2'h0; // @[LZD.scala 39:14]
  assign _T_321 = _T_319[1]; // @[LZD.scala 39:21]
  assign _T_322 = _T_319[0]; // @[LZD.scala 39:30]
  assign _T_323 = ~ _T_322; // @[LZD.scala 39:27]
  assign _T_324 = _T_321 | _T_323; // @[LZD.scala 39:25]
  assign _T_325 = {_T_320,_T_324}; // @[Cat.scala 29:58]
  assign _T_326 = _T_318[1:0]; // @[LZD.scala 44:32]
  assign _T_327 = _T_326 != 2'h0; // @[LZD.scala 39:14]
  assign _T_328 = _T_326[1]; // @[LZD.scala 39:21]
  assign _T_329 = _T_326[0]; // @[LZD.scala 39:30]
  assign _T_330 = ~ _T_329; // @[LZD.scala 39:27]
  assign _T_331 = _T_328 | _T_330; // @[LZD.scala 39:25]
  assign _T_332 = {_T_327,_T_331}; // @[Cat.scala 29:58]
  assign _T_333 = _T_325[1]; // @[Shift.scala 12:21]
  assign _T_334 = _T_332[1]; // @[Shift.scala 12:21]
  assign _T_335 = _T_333 | _T_334; // @[LZD.scala 49:16]
  assign _T_336 = ~ _T_334; // @[LZD.scala 49:27]
  assign _T_337 = _T_333 | _T_336; // @[LZD.scala 49:25]
  assign _T_338 = _T_325[0:0]; // @[LZD.scala 49:47]
  assign _T_339 = _T_332[0:0]; // @[LZD.scala 49:59]
  assign _T_340 = _T_333 ? _T_338 : _T_339; // @[LZD.scala 49:35]
  assign _T_342 = {_T_335,_T_337,_T_340}; // @[Cat.scala 29:58]
  assign _T_343 = _T_317[2]; // @[Shift.scala 12:21]
  assign _T_344 = _T_342[2]; // @[Shift.scala 12:21]
  assign _T_345 = _T_343 | _T_344; // @[LZD.scala 49:16]
  assign _T_346 = ~ _T_344; // @[LZD.scala 49:27]
  assign _T_347 = _T_343 | _T_346; // @[LZD.scala 49:25]
  assign _T_348 = _T_317[1:0]; // @[LZD.scala 49:47]
  assign _T_349 = _T_342[1:0]; // @[LZD.scala 49:59]
  assign _T_350 = _T_343 ? _T_348 : _T_349; // @[LZD.scala 49:35]
  assign _T_352 = {_T_345,_T_347,_T_350}; // @[Cat.scala 29:58]
  assign _T_353 = _T_291[7:0]; // @[LZD.scala 44:32]
  assign _T_354 = _T_353[7:4]; // @[LZD.scala 43:32]
  assign _T_355 = _T_354[3:2]; // @[LZD.scala 43:32]
  assign _T_356 = _T_355 != 2'h0; // @[LZD.scala 39:14]
  assign _T_357 = _T_355[1]; // @[LZD.scala 39:21]
  assign _T_358 = _T_355[0]; // @[LZD.scala 39:30]
  assign _T_359 = ~ _T_358; // @[LZD.scala 39:27]
  assign _T_360 = _T_357 | _T_359; // @[LZD.scala 39:25]
  assign _T_361 = {_T_356,_T_360}; // @[Cat.scala 29:58]
  assign _T_362 = _T_354[1:0]; // @[LZD.scala 44:32]
  assign _T_363 = _T_362 != 2'h0; // @[LZD.scala 39:14]
  assign _T_364 = _T_362[1]; // @[LZD.scala 39:21]
  assign _T_365 = _T_362[0]; // @[LZD.scala 39:30]
  assign _T_366 = ~ _T_365; // @[LZD.scala 39:27]
  assign _T_367 = _T_364 | _T_366; // @[LZD.scala 39:25]
  assign _T_368 = {_T_363,_T_367}; // @[Cat.scala 29:58]
  assign _T_369 = _T_361[1]; // @[Shift.scala 12:21]
  assign _T_370 = _T_368[1]; // @[Shift.scala 12:21]
  assign _T_371 = _T_369 | _T_370; // @[LZD.scala 49:16]
  assign _T_372 = ~ _T_370; // @[LZD.scala 49:27]
  assign _T_373 = _T_369 | _T_372; // @[LZD.scala 49:25]
  assign _T_374 = _T_361[0:0]; // @[LZD.scala 49:47]
  assign _T_375 = _T_368[0:0]; // @[LZD.scala 49:59]
  assign _T_376 = _T_369 ? _T_374 : _T_375; // @[LZD.scala 49:35]
  assign _T_378 = {_T_371,_T_373,_T_376}; // @[Cat.scala 29:58]
  assign _T_379 = _T_353[3:0]; // @[LZD.scala 44:32]
  assign _T_380 = _T_379[3:2]; // @[LZD.scala 43:32]
  assign _T_381 = _T_380 != 2'h0; // @[LZD.scala 39:14]
  assign _T_382 = _T_380[1]; // @[LZD.scala 39:21]
  assign _T_383 = _T_380[0]; // @[LZD.scala 39:30]
  assign _T_384 = ~ _T_383; // @[LZD.scala 39:27]
  assign _T_385 = _T_382 | _T_384; // @[LZD.scala 39:25]
  assign _T_386 = {_T_381,_T_385}; // @[Cat.scala 29:58]
  assign _T_387 = _T_379[1:0]; // @[LZD.scala 44:32]
  assign _T_388 = _T_387 != 2'h0; // @[LZD.scala 39:14]
  assign _T_389 = _T_387[1]; // @[LZD.scala 39:21]
  assign _T_390 = _T_387[0]; // @[LZD.scala 39:30]
  assign _T_391 = ~ _T_390; // @[LZD.scala 39:27]
  assign _T_392 = _T_389 | _T_391; // @[LZD.scala 39:25]
  assign _T_393 = {_T_388,_T_392}; // @[Cat.scala 29:58]
  assign _T_394 = _T_386[1]; // @[Shift.scala 12:21]
  assign _T_395 = _T_393[1]; // @[Shift.scala 12:21]
  assign _T_396 = _T_394 | _T_395; // @[LZD.scala 49:16]
  assign _T_397 = ~ _T_395; // @[LZD.scala 49:27]
  assign _T_398 = _T_394 | _T_397; // @[LZD.scala 49:25]
  assign _T_399 = _T_386[0:0]; // @[LZD.scala 49:47]
  assign _T_400 = _T_393[0:0]; // @[LZD.scala 49:59]
  assign _T_401 = _T_394 ? _T_399 : _T_400; // @[LZD.scala 49:35]
  assign _T_403 = {_T_396,_T_398,_T_401}; // @[Cat.scala 29:58]
  assign _T_404 = _T_378[2]; // @[Shift.scala 12:21]
  assign _T_405 = _T_403[2]; // @[Shift.scala 12:21]
  assign _T_406 = _T_404 | _T_405; // @[LZD.scala 49:16]
  assign _T_407 = ~ _T_405; // @[LZD.scala 49:27]
  assign _T_408 = _T_404 | _T_407; // @[LZD.scala 49:25]
  assign _T_409 = _T_378[1:0]; // @[LZD.scala 49:47]
  assign _T_410 = _T_403[1:0]; // @[LZD.scala 49:59]
  assign _T_411 = _T_404 ? _T_409 : _T_410; // @[LZD.scala 49:35]
  assign _T_413 = {_T_406,_T_408,_T_411}; // @[Cat.scala 29:58]
  assign _T_414 = _T_352[3]; // @[Shift.scala 12:21]
  assign _T_415 = _T_413[3]; // @[Shift.scala 12:21]
  assign _T_416 = _T_414 | _T_415; // @[LZD.scala 49:16]
  assign _T_417 = ~ _T_415; // @[LZD.scala 49:27]
  assign _T_418 = _T_414 | _T_417; // @[LZD.scala 49:25]
  assign _T_419 = _T_352[2:0]; // @[LZD.scala 49:47]
  assign _T_420 = _T_413[2:0]; // @[LZD.scala 49:59]
  assign _T_421 = _T_414 ? _T_419 : _T_420; // @[LZD.scala 49:35]
  assign _T_423 = {_T_416,_T_418,_T_421}; // @[Cat.scala 29:58]
  assign _T_424 = _T_290[15:0]; // @[LZD.scala 44:32]
  assign _T_425 = _T_424[15:8]; // @[LZD.scala 43:32]
  assign _T_426 = _T_425[7:4]; // @[LZD.scala 43:32]
  assign _T_427 = _T_426[3:2]; // @[LZD.scala 43:32]
  assign _T_428 = _T_427 != 2'h0; // @[LZD.scala 39:14]
  assign _T_429 = _T_427[1]; // @[LZD.scala 39:21]
  assign _T_430 = _T_427[0]; // @[LZD.scala 39:30]
  assign _T_431 = ~ _T_430; // @[LZD.scala 39:27]
  assign _T_432 = _T_429 | _T_431; // @[LZD.scala 39:25]
  assign _T_433 = {_T_428,_T_432}; // @[Cat.scala 29:58]
  assign _T_434 = _T_426[1:0]; // @[LZD.scala 44:32]
  assign _T_435 = _T_434 != 2'h0; // @[LZD.scala 39:14]
  assign _T_436 = _T_434[1]; // @[LZD.scala 39:21]
  assign _T_437 = _T_434[0]; // @[LZD.scala 39:30]
  assign _T_438 = ~ _T_437; // @[LZD.scala 39:27]
  assign _T_439 = _T_436 | _T_438; // @[LZD.scala 39:25]
  assign _T_440 = {_T_435,_T_439}; // @[Cat.scala 29:58]
  assign _T_441 = _T_433[1]; // @[Shift.scala 12:21]
  assign _T_442 = _T_440[1]; // @[Shift.scala 12:21]
  assign _T_443 = _T_441 | _T_442; // @[LZD.scala 49:16]
  assign _T_444 = ~ _T_442; // @[LZD.scala 49:27]
  assign _T_445 = _T_441 | _T_444; // @[LZD.scala 49:25]
  assign _T_446 = _T_433[0:0]; // @[LZD.scala 49:47]
  assign _T_447 = _T_440[0:0]; // @[LZD.scala 49:59]
  assign _T_448 = _T_441 ? _T_446 : _T_447; // @[LZD.scala 49:35]
  assign _T_450 = {_T_443,_T_445,_T_448}; // @[Cat.scala 29:58]
  assign _T_451 = _T_425[3:0]; // @[LZD.scala 44:32]
  assign _T_452 = _T_451[3:2]; // @[LZD.scala 43:32]
  assign _T_453 = _T_452 != 2'h0; // @[LZD.scala 39:14]
  assign _T_454 = _T_452[1]; // @[LZD.scala 39:21]
  assign _T_455 = _T_452[0]; // @[LZD.scala 39:30]
  assign _T_456 = ~ _T_455; // @[LZD.scala 39:27]
  assign _T_457 = _T_454 | _T_456; // @[LZD.scala 39:25]
  assign _T_458 = {_T_453,_T_457}; // @[Cat.scala 29:58]
  assign _T_459 = _T_451[1:0]; // @[LZD.scala 44:32]
  assign _T_460 = _T_459 != 2'h0; // @[LZD.scala 39:14]
  assign _T_461 = _T_459[1]; // @[LZD.scala 39:21]
  assign _T_462 = _T_459[0]; // @[LZD.scala 39:30]
  assign _T_463 = ~ _T_462; // @[LZD.scala 39:27]
  assign _T_464 = _T_461 | _T_463; // @[LZD.scala 39:25]
  assign _T_465 = {_T_460,_T_464}; // @[Cat.scala 29:58]
  assign _T_466 = _T_458[1]; // @[Shift.scala 12:21]
  assign _T_467 = _T_465[1]; // @[Shift.scala 12:21]
  assign _T_468 = _T_466 | _T_467; // @[LZD.scala 49:16]
  assign _T_469 = ~ _T_467; // @[LZD.scala 49:27]
  assign _T_470 = _T_466 | _T_469; // @[LZD.scala 49:25]
  assign _T_471 = _T_458[0:0]; // @[LZD.scala 49:47]
  assign _T_472 = _T_465[0:0]; // @[LZD.scala 49:59]
  assign _T_473 = _T_466 ? _T_471 : _T_472; // @[LZD.scala 49:35]
  assign _T_475 = {_T_468,_T_470,_T_473}; // @[Cat.scala 29:58]
  assign _T_476 = _T_450[2]; // @[Shift.scala 12:21]
  assign _T_477 = _T_475[2]; // @[Shift.scala 12:21]
  assign _T_478 = _T_476 | _T_477; // @[LZD.scala 49:16]
  assign _T_479 = ~ _T_477; // @[LZD.scala 49:27]
  assign _T_480 = _T_476 | _T_479; // @[LZD.scala 49:25]
  assign _T_481 = _T_450[1:0]; // @[LZD.scala 49:47]
  assign _T_482 = _T_475[1:0]; // @[LZD.scala 49:59]
  assign _T_483 = _T_476 ? _T_481 : _T_482; // @[LZD.scala 49:35]
  assign _T_485 = {_T_478,_T_480,_T_483}; // @[Cat.scala 29:58]
  assign _T_486 = _T_424[7:0]; // @[LZD.scala 44:32]
  assign _T_487 = _T_486[7:4]; // @[LZD.scala 43:32]
  assign _T_488 = _T_487[3:2]; // @[LZD.scala 43:32]
  assign _T_489 = _T_488 != 2'h0; // @[LZD.scala 39:14]
  assign _T_490 = _T_488[1]; // @[LZD.scala 39:21]
  assign _T_491 = _T_488[0]; // @[LZD.scala 39:30]
  assign _T_492 = ~ _T_491; // @[LZD.scala 39:27]
  assign _T_493 = _T_490 | _T_492; // @[LZD.scala 39:25]
  assign _T_494 = {_T_489,_T_493}; // @[Cat.scala 29:58]
  assign _T_495 = _T_487[1:0]; // @[LZD.scala 44:32]
  assign _T_496 = _T_495 != 2'h0; // @[LZD.scala 39:14]
  assign _T_497 = _T_495[1]; // @[LZD.scala 39:21]
  assign _T_498 = _T_495[0]; // @[LZD.scala 39:30]
  assign _T_499 = ~ _T_498; // @[LZD.scala 39:27]
  assign _T_500 = _T_497 | _T_499; // @[LZD.scala 39:25]
  assign _T_501 = {_T_496,_T_500}; // @[Cat.scala 29:58]
  assign _T_502 = _T_494[1]; // @[Shift.scala 12:21]
  assign _T_503 = _T_501[1]; // @[Shift.scala 12:21]
  assign _T_504 = _T_502 | _T_503; // @[LZD.scala 49:16]
  assign _T_505 = ~ _T_503; // @[LZD.scala 49:27]
  assign _T_506 = _T_502 | _T_505; // @[LZD.scala 49:25]
  assign _T_507 = _T_494[0:0]; // @[LZD.scala 49:47]
  assign _T_508 = _T_501[0:0]; // @[LZD.scala 49:59]
  assign _T_509 = _T_502 ? _T_507 : _T_508; // @[LZD.scala 49:35]
  assign _T_511 = {_T_504,_T_506,_T_509}; // @[Cat.scala 29:58]
  assign _T_512 = _T_486[3:0]; // @[LZD.scala 44:32]
  assign _T_513 = _T_512[3:2]; // @[LZD.scala 43:32]
  assign _T_514 = _T_513 != 2'h0; // @[LZD.scala 39:14]
  assign _T_515 = _T_513[1]; // @[LZD.scala 39:21]
  assign _T_516 = _T_513[0]; // @[LZD.scala 39:30]
  assign _T_517 = ~ _T_516; // @[LZD.scala 39:27]
  assign _T_518 = _T_515 | _T_517; // @[LZD.scala 39:25]
  assign _T_519 = {_T_514,_T_518}; // @[Cat.scala 29:58]
  assign _T_520 = _T_512[1:0]; // @[LZD.scala 44:32]
  assign _T_521 = _T_520 != 2'h0; // @[LZD.scala 39:14]
  assign _T_522 = _T_520[1]; // @[LZD.scala 39:21]
  assign _T_523 = _T_520[0]; // @[LZD.scala 39:30]
  assign _T_524 = ~ _T_523; // @[LZD.scala 39:27]
  assign _T_525 = _T_522 | _T_524; // @[LZD.scala 39:25]
  assign _T_526 = {_T_521,_T_525}; // @[Cat.scala 29:58]
  assign _T_527 = _T_519[1]; // @[Shift.scala 12:21]
  assign _T_528 = _T_526[1]; // @[Shift.scala 12:21]
  assign _T_529 = _T_527 | _T_528; // @[LZD.scala 49:16]
  assign _T_530 = ~ _T_528; // @[LZD.scala 49:27]
  assign _T_531 = _T_527 | _T_530; // @[LZD.scala 49:25]
  assign _T_532 = _T_519[0:0]; // @[LZD.scala 49:47]
  assign _T_533 = _T_526[0:0]; // @[LZD.scala 49:59]
  assign _T_534 = _T_527 ? _T_532 : _T_533; // @[LZD.scala 49:35]
  assign _T_536 = {_T_529,_T_531,_T_534}; // @[Cat.scala 29:58]
  assign _T_537 = _T_511[2]; // @[Shift.scala 12:21]
  assign _T_538 = _T_536[2]; // @[Shift.scala 12:21]
  assign _T_539 = _T_537 | _T_538; // @[LZD.scala 49:16]
  assign _T_540 = ~ _T_538; // @[LZD.scala 49:27]
  assign _T_541 = _T_537 | _T_540; // @[LZD.scala 49:25]
  assign _T_542 = _T_511[1:0]; // @[LZD.scala 49:47]
  assign _T_543 = _T_536[1:0]; // @[LZD.scala 49:59]
  assign _T_544 = _T_537 ? _T_542 : _T_543; // @[LZD.scala 49:35]
  assign _T_546 = {_T_539,_T_541,_T_544}; // @[Cat.scala 29:58]
  assign _T_547 = _T_485[3]; // @[Shift.scala 12:21]
  assign _T_548 = _T_546[3]; // @[Shift.scala 12:21]
  assign _T_549 = _T_547 | _T_548; // @[LZD.scala 49:16]
  assign _T_550 = ~ _T_548; // @[LZD.scala 49:27]
  assign _T_551 = _T_547 | _T_550; // @[LZD.scala 49:25]
  assign _T_552 = _T_485[2:0]; // @[LZD.scala 49:47]
  assign _T_553 = _T_546[2:0]; // @[LZD.scala 49:59]
  assign _T_554 = _T_547 ? _T_552 : _T_553; // @[LZD.scala 49:35]
  assign _T_556 = {_T_549,_T_551,_T_554}; // @[Cat.scala 29:58]
  assign _T_557 = _T_423[4]; // @[Shift.scala 12:21]
  assign _T_558 = _T_556[4]; // @[Shift.scala 12:21]
  assign _T_559 = _T_557 | _T_558; // @[LZD.scala 49:16]
  assign _T_560 = ~ _T_558; // @[LZD.scala 49:27]
  assign _T_561 = _T_557 | _T_560; // @[LZD.scala 49:25]
  assign _T_562 = _T_423[3:0]; // @[LZD.scala 49:47]
  assign _T_563 = _T_556[3:0]; // @[LZD.scala 49:59]
  assign _T_564 = _T_557 ? _T_562 : _T_563; // @[LZD.scala 49:35]
  assign _T_566 = {_T_559,_T_561,_T_564}; // @[Cat.scala 29:58]
  assign _T_567 = _T_289[5]; // @[Shift.scala 12:21]
  assign _T_568 = _T_566[5]; // @[Shift.scala 12:21]
  assign _T_569 = _T_567 | _T_568; // @[LZD.scala 49:16]
  assign _T_570 = ~ _T_568; // @[LZD.scala 49:27]
  assign _T_571 = _T_567 | _T_570; // @[LZD.scala 49:25]
  assign _T_572 = _T_289[4:0]; // @[LZD.scala 49:47]
  assign _T_573 = _T_566[4:0]; // @[LZD.scala 49:59]
  assign _T_574 = _T_567 ? _T_572 : _T_573; // @[LZD.scala 49:35]
  assign _T_576 = {_T_569,_T_571,_T_574}; // @[Cat.scala 29:58]
  assign _T_577 = _T_11[63:0]; // @[LZD.scala 44:32]
  assign _T_578 = _T_577[63:32]; // @[LZD.scala 43:32]
  assign _T_579 = _T_578[31:16]; // @[LZD.scala 43:32]
  assign _T_580 = _T_579[15:8]; // @[LZD.scala 43:32]
  assign _T_581 = _T_580[7:4]; // @[LZD.scala 43:32]
  assign _T_582 = _T_581[3:2]; // @[LZD.scala 43:32]
  assign _T_583 = _T_582 != 2'h0; // @[LZD.scala 39:14]
  assign _T_584 = _T_582[1]; // @[LZD.scala 39:21]
  assign _T_585 = _T_582[0]; // @[LZD.scala 39:30]
  assign _T_586 = ~ _T_585; // @[LZD.scala 39:27]
  assign _T_587 = _T_584 | _T_586; // @[LZD.scala 39:25]
  assign _T_588 = {_T_583,_T_587}; // @[Cat.scala 29:58]
  assign _T_589 = _T_581[1:0]; // @[LZD.scala 44:32]
  assign _T_590 = _T_589 != 2'h0; // @[LZD.scala 39:14]
  assign _T_591 = _T_589[1]; // @[LZD.scala 39:21]
  assign _T_592 = _T_589[0]; // @[LZD.scala 39:30]
  assign _T_593 = ~ _T_592; // @[LZD.scala 39:27]
  assign _T_594 = _T_591 | _T_593; // @[LZD.scala 39:25]
  assign _T_595 = {_T_590,_T_594}; // @[Cat.scala 29:58]
  assign _T_596 = _T_588[1]; // @[Shift.scala 12:21]
  assign _T_597 = _T_595[1]; // @[Shift.scala 12:21]
  assign _T_598 = _T_596 | _T_597; // @[LZD.scala 49:16]
  assign _T_599 = ~ _T_597; // @[LZD.scala 49:27]
  assign _T_600 = _T_596 | _T_599; // @[LZD.scala 49:25]
  assign _T_601 = _T_588[0:0]; // @[LZD.scala 49:47]
  assign _T_602 = _T_595[0:0]; // @[LZD.scala 49:59]
  assign _T_603 = _T_596 ? _T_601 : _T_602; // @[LZD.scala 49:35]
  assign _T_605 = {_T_598,_T_600,_T_603}; // @[Cat.scala 29:58]
  assign _T_606 = _T_580[3:0]; // @[LZD.scala 44:32]
  assign _T_607 = _T_606[3:2]; // @[LZD.scala 43:32]
  assign _T_608 = _T_607 != 2'h0; // @[LZD.scala 39:14]
  assign _T_609 = _T_607[1]; // @[LZD.scala 39:21]
  assign _T_610 = _T_607[0]; // @[LZD.scala 39:30]
  assign _T_611 = ~ _T_610; // @[LZD.scala 39:27]
  assign _T_612 = _T_609 | _T_611; // @[LZD.scala 39:25]
  assign _T_613 = {_T_608,_T_612}; // @[Cat.scala 29:58]
  assign _T_614 = _T_606[1:0]; // @[LZD.scala 44:32]
  assign _T_615 = _T_614 != 2'h0; // @[LZD.scala 39:14]
  assign _T_616 = _T_614[1]; // @[LZD.scala 39:21]
  assign _T_617 = _T_614[0]; // @[LZD.scala 39:30]
  assign _T_618 = ~ _T_617; // @[LZD.scala 39:27]
  assign _T_619 = _T_616 | _T_618; // @[LZD.scala 39:25]
  assign _T_620 = {_T_615,_T_619}; // @[Cat.scala 29:58]
  assign _T_621 = _T_613[1]; // @[Shift.scala 12:21]
  assign _T_622 = _T_620[1]; // @[Shift.scala 12:21]
  assign _T_623 = _T_621 | _T_622; // @[LZD.scala 49:16]
  assign _T_624 = ~ _T_622; // @[LZD.scala 49:27]
  assign _T_625 = _T_621 | _T_624; // @[LZD.scala 49:25]
  assign _T_626 = _T_613[0:0]; // @[LZD.scala 49:47]
  assign _T_627 = _T_620[0:0]; // @[LZD.scala 49:59]
  assign _T_628 = _T_621 ? _T_626 : _T_627; // @[LZD.scala 49:35]
  assign _T_630 = {_T_623,_T_625,_T_628}; // @[Cat.scala 29:58]
  assign _T_631 = _T_605[2]; // @[Shift.scala 12:21]
  assign _T_632 = _T_630[2]; // @[Shift.scala 12:21]
  assign _T_633 = _T_631 | _T_632; // @[LZD.scala 49:16]
  assign _T_634 = ~ _T_632; // @[LZD.scala 49:27]
  assign _T_635 = _T_631 | _T_634; // @[LZD.scala 49:25]
  assign _T_636 = _T_605[1:0]; // @[LZD.scala 49:47]
  assign _T_637 = _T_630[1:0]; // @[LZD.scala 49:59]
  assign _T_638 = _T_631 ? _T_636 : _T_637; // @[LZD.scala 49:35]
  assign _T_640 = {_T_633,_T_635,_T_638}; // @[Cat.scala 29:58]
  assign _T_641 = _T_579[7:0]; // @[LZD.scala 44:32]
  assign _T_642 = _T_641[7:4]; // @[LZD.scala 43:32]
  assign _T_643 = _T_642[3:2]; // @[LZD.scala 43:32]
  assign _T_644 = _T_643 != 2'h0; // @[LZD.scala 39:14]
  assign _T_645 = _T_643[1]; // @[LZD.scala 39:21]
  assign _T_646 = _T_643[0]; // @[LZD.scala 39:30]
  assign _T_647 = ~ _T_646; // @[LZD.scala 39:27]
  assign _T_648 = _T_645 | _T_647; // @[LZD.scala 39:25]
  assign _T_649 = {_T_644,_T_648}; // @[Cat.scala 29:58]
  assign _T_650 = _T_642[1:0]; // @[LZD.scala 44:32]
  assign _T_651 = _T_650 != 2'h0; // @[LZD.scala 39:14]
  assign _T_652 = _T_650[1]; // @[LZD.scala 39:21]
  assign _T_653 = _T_650[0]; // @[LZD.scala 39:30]
  assign _T_654 = ~ _T_653; // @[LZD.scala 39:27]
  assign _T_655 = _T_652 | _T_654; // @[LZD.scala 39:25]
  assign _T_656 = {_T_651,_T_655}; // @[Cat.scala 29:58]
  assign _T_657 = _T_649[1]; // @[Shift.scala 12:21]
  assign _T_658 = _T_656[1]; // @[Shift.scala 12:21]
  assign _T_659 = _T_657 | _T_658; // @[LZD.scala 49:16]
  assign _T_660 = ~ _T_658; // @[LZD.scala 49:27]
  assign _T_661 = _T_657 | _T_660; // @[LZD.scala 49:25]
  assign _T_662 = _T_649[0:0]; // @[LZD.scala 49:47]
  assign _T_663 = _T_656[0:0]; // @[LZD.scala 49:59]
  assign _T_664 = _T_657 ? _T_662 : _T_663; // @[LZD.scala 49:35]
  assign _T_666 = {_T_659,_T_661,_T_664}; // @[Cat.scala 29:58]
  assign _T_667 = _T_641[3:0]; // @[LZD.scala 44:32]
  assign _T_668 = _T_667[3:2]; // @[LZD.scala 43:32]
  assign _T_669 = _T_668 != 2'h0; // @[LZD.scala 39:14]
  assign _T_670 = _T_668[1]; // @[LZD.scala 39:21]
  assign _T_671 = _T_668[0]; // @[LZD.scala 39:30]
  assign _T_672 = ~ _T_671; // @[LZD.scala 39:27]
  assign _T_673 = _T_670 | _T_672; // @[LZD.scala 39:25]
  assign _T_674 = {_T_669,_T_673}; // @[Cat.scala 29:58]
  assign _T_675 = _T_667[1:0]; // @[LZD.scala 44:32]
  assign _T_676 = _T_675 != 2'h0; // @[LZD.scala 39:14]
  assign _T_677 = _T_675[1]; // @[LZD.scala 39:21]
  assign _T_678 = _T_675[0]; // @[LZD.scala 39:30]
  assign _T_679 = ~ _T_678; // @[LZD.scala 39:27]
  assign _T_680 = _T_677 | _T_679; // @[LZD.scala 39:25]
  assign _T_681 = {_T_676,_T_680}; // @[Cat.scala 29:58]
  assign _T_682 = _T_674[1]; // @[Shift.scala 12:21]
  assign _T_683 = _T_681[1]; // @[Shift.scala 12:21]
  assign _T_684 = _T_682 | _T_683; // @[LZD.scala 49:16]
  assign _T_685 = ~ _T_683; // @[LZD.scala 49:27]
  assign _T_686 = _T_682 | _T_685; // @[LZD.scala 49:25]
  assign _T_687 = _T_674[0:0]; // @[LZD.scala 49:47]
  assign _T_688 = _T_681[0:0]; // @[LZD.scala 49:59]
  assign _T_689 = _T_682 ? _T_687 : _T_688; // @[LZD.scala 49:35]
  assign _T_691 = {_T_684,_T_686,_T_689}; // @[Cat.scala 29:58]
  assign _T_692 = _T_666[2]; // @[Shift.scala 12:21]
  assign _T_693 = _T_691[2]; // @[Shift.scala 12:21]
  assign _T_694 = _T_692 | _T_693; // @[LZD.scala 49:16]
  assign _T_695 = ~ _T_693; // @[LZD.scala 49:27]
  assign _T_696 = _T_692 | _T_695; // @[LZD.scala 49:25]
  assign _T_697 = _T_666[1:0]; // @[LZD.scala 49:47]
  assign _T_698 = _T_691[1:0]; // @[LZD.scala 49:59]
  assign _T_699 = _T_692 ? _T_697 : _T_698; // @[LZD.scala 49:35]
  assign _T_701 = {_T_694,_T_696,_T_699}; // @[Cat.scala 29:58]
  assign _T_702 = _T_640[3]; // @[Shift.scala 12:21]
  assign _T_703 = _T_701[3]; // @[Shift.scala 12:21]
  assign _T_704 = _T_702 | _T_703; // @[LZD.scala 49:16]
  assign _T_705 = ~ _T_703; // @[LZD.scala 49:27]
  assign _T_706 = _T_702 | _T_705; // @[LZD.scala 49:25]
  assign _T_707 = _T_640[2:0]; // @[LZD.scala 49:47]
  assign _T_708 = _T_701[2:0]; // @[LZD.scala 49:59]
  assign _T_709 = _T_702 ? _T_707 : _T_708; // @[LZD.scala 49:35]
  assign _T_711 = {_T_704,_T_706,_T_709}; // @[Cat.scala 29:58]
  assign _T_712 = _T_578[15:0]; // @[LZD.scala 44:32]
  assign _T_713 = _T_712[15:8]; // @[LZD.scala 43:32]
  assign _T_714 = _T_713[7:4]; // @[LZD.scala 43:32]
  assign _T_715 = _T_714[3:2]; // @[LZD.scala 43:32]
  assign _T_716 = _T_715 != 2'h0; // @[LZD.scala 39:14]
  assign _T_717 = _T_715[1]; // @[LZD.scala 39:21]
  assign _T_718 = _T_715[0]; // @[LZD.scala 39:30]
  assign _T_719 = ~ _T_718; // @[LZD.scala 39:27]
  assign _T_720 = _T_717 | _T_719; // @[LZD.scala 39:25]
  assign _T_721 = {_T_716,_T_720}; // @[Cat.scala 29:58]
  assign _T_722 = _T_714[1:0]; // @[LZD.scala 44:32]
  assign _T_723 = _T_722 != 2'h0; // @[LZD.scala 39:14]
  assign _T_724 = _T_722[1]; // @[LZD.scala 39:21]
  assign _T_725 = _T_722[0]; // @[LZD.scala 39:30]
  assign _T_726 = ~ _T_725; // @[LZD.scala 39:27]
  assign _T_727 = _T_724 | _T_726; // @[LZD.scala 39:25]
  assign _T_728 = {_T_723,_T_727}; // @[Cat.scala 29:58]
  assign _T_729 = _T_721[1]; // @[Shift.scala 12:21]
  assign _T_730 = _T_728[1]; // @[Shift.scala 12:21]
  assign _T_731 = _T_729 | _T_730; // @[LZD.scala 49:16]
  assign _T_732 = ~ _T_730; // @[LZD.scala 49:27]
  assign _T_733 = _T_729 | _T_732; // @[LZD.scala 49:25]
  assign _T_734 = _T_721[0:0]; // @[LZD.scala 49:47]
  assign _T_735 = _T_728[0:0]; // @[LZD.scala 49:59]
  assign _T_736 = _T_729 ? _T_734 : _T_735; // @[LZD.scala 49:35]
  assign _T_738 = {_T_731,_T_733,_T_736}; // @[Cat.scala 29:58]
  assign _T_739 = _T_713[3:0]; // @[LZD.scala 44:32]
  assign _T_740 = _T_739[3:2]; // @[LZD.scala 43:32]
  assign _T_741 = _T_740 != 2'h0; // @[LZD.scala 39:14]
  assign _T_742 = _T_740[1]; // @[LZD.scala 39:21]
  assign _T_743 = _T_740[0]; // @[LZD.scala 39:30]
  assign _T_744 = ~ _T_743; // @[LZD.scala 39:27]
  assign _T_745 = _T_742 | _T_744; // @[LZD.scala 39:25]
  assign _T_746 = {_T_741,_T_745}; // @[Cat.scala 29:58]
  assign _T_747 = _T_739[1:0]; // @[LZD.scala 44:32]
  assign _T_748 = _T_747 != 2'h0; // @[LZD.scala 39:14]
  assign _T_749 = _T_747[1]; // @[LZD.scala 39:21]
  assign _T_750 = _T_747[0]; // @[LZD.scala 39:30]
  assign _T_751 = ~ _T_750; // @[LZD.scala 39:27]
  assign _T_752 = _T_749 | _T_751; // @[LZD.scala 39:25]
  assign _T_753 = {_T_748,_T_752}; // @[Cat.scala 29:58]
  assign _T_754 = _T_746[1]; // @[Shift.scala 12:21]
  assign _T_755 = _T_753[1]; // @[Shift.scala 12:21]
  assign _T_756 = _T_754 | _T_755; // @[LZD.scala 49:16]
  assign _T_757 = ~ _T_755; // @[LZD.scala 49:27]
  assign _T_758 = _T_754 | _T_757; // @[LZD.scala 49:25]
  assign _T_759 = _T_746[0:0]; // @[LZD.scala 49:47]
  assign _T_760 = _T_753[0:0]; // @[LZD.scala 49:59]
  assign _T_761 = _T_754 ? _T_759 : _T_760; // @[LZD.scala 49:35]
  assign _T_763 = {_T_756,_T_758,_T_761}; // @[Cat.scala 29:58]
  assign _T_764 = _T_738[2]; // @[Shift.scala 12:21]
  assign _T_765 = _T_763[2]; // @[Shift.scala 12:21]
  assign _T_766 = _T_764 | _T_765; // @[LZD.scala 49:16]
  assign _T_767 = ~ _T_765; // @[LZD.scala 49:27]
  assign _T_768 = _T_764 | _T_767; // @[LZD.scala 49:25]
  assign _T_769 = _T_738[1:0]; // @[LZD.scala 49:47]
  assign _T_770 = _T_763[1:0]; // @[LZD.scala 49:59]
  assign _T_771 = _T_764 ? _T_769 : _T_770; // @[LZD.scala 49:35]
  assign _T_773 = {_T_766,_T_768,_T_771}; // @[Cat.scala 29:58]
  assign _T_774 = _T_712[7:0]; // @[LZD.scala 44:32]
  assign _T_775 = _T_774[7:4]; // @[LZD.scala 43:32]
  assign _T_776 = _T_775[3:2]; // @[LZD.scala 43:32]
  assign _T_777 = _T_776 != 2'h0; // @[LZD.scala 39:14]
  assign _T_778 = _T_776[1]; // @[LZD.scala 39:21]
  assign _T_779 = _T_776[0]; // @[LZD.scala 39:30]
  assign _T_780 = ~ _T_779; // @[LZD.scala 39:27]
  assign _T_781 = _T_778 | _T_780; // @[LZD.scala 39:25]
  assign _T_782 = {_T_777,_T_781}; // @[Cat.scala 29:58]
  assign _T_783 = _T_775[1:0]; // @[LZD.scala 44:32]
  assign _T_784 = _T_783 != 2'h0; // @[LZD.scala 39:14]
  assign _T_785 = _T_783[1]; // @[LZD.scala 39:21]
  assign _T_786 = _T_783[0]; // @[LZD.scala 39:30]
  assign _T_787 = ~ _T_786; // @[LZD.scala 39:27]
  assign _T_788 = _T_785 | _T_787; // @[LZD.scala 39:25]
  assign _T_789 = {_T_784,_T_788}; // @[Cat.scala 29:58]
  assign _T_790 = _T_782[1]; // @[Shift.scala 12:21]
  assign _T_791 = _T_789[1]; // @[Shift.scala 12:21]
  assign _T_792 = _T_790 | _T_791; // @[LZD.scala 49:16]
  assign _T_793 = ~ _T_791; // @[LZD.scala 49:27]
  assign _T_794 = _T_790 | _T_793; // @[LZD.scala 49:25]
  assign _T_795 = _T_782[0:0]; // @[LZD.scala 49:47]
  assign _T_796 = _T_789[0:0]; // @[LZD.scala 49:59]
  assign _T_797 = _T_790 ? _T_795 : _T_796; // @[LZD.scala 49:35]
  assign _T_799 = {_T_792,_T_794,_T_797}; // @[Cat.scala 29:58]
  assign _T_800 = _T_774[3:0]; // @[LZD.scala 44:32]
  assign _T_801 = _T_800[3:2]; // @[LZD.scala 43:32]
  assign _T_802 = _T_801 != 2'h0; // @[LZD.scala 39:14]
  assign _T_803 = _T_801[1]; // @[LZD.scala 39:21]
  assign _T_804 = _T_801[0]; // @[LZD.scala 39:30]
  assign _T_805 = ~ _T_804; // @[LZD.scala 39:27]
  assign _T_806 = _T_803 | _T_805; // @[LZD.scala 39:25]
  assign _T_807 = {_T_802,_T_806}; // @[Cat.scala 29:58]
  assign _T_808 = _T_800[1:0]; // @[LZD.scala 44:32]
  assign _T_809 = _T_808 != 2'h0; // @[LZD.scala 39:14]
  assign _T_810 = _T_808[1]; // @[LZD.scala 39:21]
  assign _T_811 = _T_808[0]; // @[LZD.scala 39:30]
  assign _T_812 = ~ _T_811; // @[LZD.scala 39:27]
  assign _T_813 = _T_810 | _T_812; // @[LZD.scala 39:25]
  assign _T_814 = {_T_809,_T_813}; // @[Cat.scala 29:58]
  assign _T_815 = _T_807[1]; // @[Shift.scala 12:21]
  assign _T_816 = _T_814[1]; // @[Shift.scala 12:21]
  assign _T_817 = _T_815 | _T_816; // @[LZD.scala 49:16]
  assign _T_818 = ~ _T_816; // @[LZD.scala 49:27]
  assign _T_819 = _T_815 | _T_818; // @[LZD.scala 49:25]
  assign _T_820 = _T_807[0:0]; // @[LZD.scala 49:47]
  assign _T_821 = _T_814[0:0]; // @[LZD.scala 49:59]
  assign _T_822 = _T_815 ? _T_820 : _T_821; // @[LZD.scala 49:35]
  assign _T_824 = {_T_817,_T_819,_T_822}; // @[Cat.scala 29:58]
  assign _T_825 = _T_799[2]; // @[Shift.scala 12:21]
  assign _T_826 = _T_824[2]; // @[Shift.scala 12:21]
  assign _T_827 = _T_825 | _T_826; // @[LZD.scala 49:16]
  assign _T_828 = ~ _T_826; // @[LZD.scala 49:27]
  assign _T_829 = _T_825 | _T_828; // @[LZD.scala 49:25]
  assign _T_830 = _T_799[1:0]; // @[LZD.scala 49:47]
  assign _T_831 = _T_824[1:0]; // @[LZD.scala 49:59]
  assign _T_832 = _T_825 ? _T_830 : _T_831; // @[LZD.scala 49:35]
  assign _T_834 = {_T_827,_T_829,_T_832}; // @[Cat.scala 29:58]
  assign _T_835 = _T_773[3]; // @[Shift.scala 12:21]
  assign _T_836 = _T_834[3]; // @[Shift.scala 12:21]
  assign _T_837 = _T_835 | _T_836; // @[LZD.scala 49:16]
  assign _T_838 = ~ _T_836; // @[LZD.scala 49:27]
  assign _T_839 = _T_835 | _T_838; // @[LZD.scala 49:25]
  assign _T_840 = _T_773[2:0]; // @[LZD.scala 49:47]
  assign _T_841 = _T_834[2:0]; // @[LZD.scala 49:59]
  assign _T_842 = _T_835 ? _T_840 : _T_841; // @[LZD.scala 49:35]
  assign _T_844 = {_T_837,_T_839,_T_842}; // @[Cat.scala 29:58]
  assign _T_845 = _T_711[4]; // @[Shift.scala 12:21]
  assign _T_846 = _T_844[4]; // @[Shift.scala 12:21]
  assign _T_847 = _T_845 | _T_846; // @[LZD.scala 49:16]
  assign _T_848 = ~ _T_846; // @[LZD.scala 49:27]
  assign _T_849 = _T_845 | _T_848; // @[LZD.scala 49:25]
  assign _T_850 = _T_711[3:0]; // @[LZD.scala 49:47]
  assign _T_851 = _T_844[3:0]; // @[LZD.scala 49:59]
  assign _T_852 = _T_845 ? _T_850 : _T_851; // @[LZD.scala 49:35]
  assign _T_854 = {_T_847,_T_849,_T_852}; // @[Cat.scala 29:58]
  assign _T_855 = _T_577[31:0]; // @[LZD.scala 44:32]
  assign _T_856 = _T_855[31:16]; // @[LZD.scala 43:32]
  assign _T_857 = _T_856[15:8]; // @[LZD.scala 43:32]
  assign _T_858 = _T_857[7:4]; // @[LZD.scala 43:32]
  assign _T_859 = _T_858[3:2]; // @[LZD.scala 43:32]
  assign _T_860 = _T_859 != 2'h0; // @[LZD.scala 39:14]
  assign _T_861 = _T_859[1]; // @[LZD.scala 39:21]
  assign _T_862 = _T_859[0]; // @[LZD.scala 39:30]
  assign _T_863 = ~ _T_862; // @[LZD.scala 39:27]
  assign _T_864 = _T_861 | _T_863; // @[LZD.scala 39:25]
  assign _T_865 = {_T_860,_T_864}; // @[Cat.scala 29:58]
  assign _T_866 = _T_858[1:0]; // @[LZD.scala 44:32]
  assign _T_867 = _T_866 != 2'h0; // @[LZD.scala 39:14]
  assign _T_868 = _T_866[1]; // @[LZD.scala 39:21]
  assign _T_869 = _T_866[0]; // @[LZD.scala 39:30]
  assign _T_870 = ~ _T_869; // @[LZD.scala 39:27]
  assign _T_871 = _T_868 | _T_870; // @[LZD.scala 39:25]
  assign _T_872 = {_T_867,_T_871}; // @[Cat.scala 29:58]
  assign _T_873 = _T_865[1]; // @[Shift.scala 12:21]
  assign _T_874 = _T_872[1]; // @[Shift.scala 12:21]
  assign _T_875 = _T_873 | _T_874; // @[LZD.scala 49:16]
  assign _T_876 = ~ _T_874; // @[LZD.scala 49:27]
  assign _T_877 = _T_873 | _T_876; // @[LZD.scala 49:25]
  assign _T_878 = _T_865[0:0]; // @[LZD.scala 49:47]
  assign _T_879 = _T_872[0:0]; // @[LZD.scala 49:59]
  assign _T_880 = _T_873 ? _T_878 : _T_879; // @[LZD.scala 49:35]
  assign _T_882 = {_T_875,_T_877,_T_880}; // @[Cat.scala 29:58]
  assign _T_883 = _T_857[3:0]; // @[LZD.scala 44:32]
  assign _T_884 = _T_883[3:2]; // @[LZD.scala 43:32]
  assign _T_885 = _T_884 != 2'h0; // @[LZD.scala 39:14]
  assign _T_886 = _T_884[1]; // @[LZD.scala 39:21]
  assign _T_887 = _T_884[0]; // @[LZD.scala 39:30]
  assign _T_888 = ~ _T_887; // @[LZD.scala 39:27]
  assign _T_889 = _T_886 | _T_888; // @[LZD.scala 39:25]
  assign _T_890 = {_T_885,_T_889}; // @[Cat.scala 29:58]
  assign _T_891 = _T_883[1:0]; // @[LZD.scala 44:32]
  assign _T_892 = _T_891 != 2'h0; // @[LZD.scala 39:14]
  assign _T_893 = _T_891[1]; // @[LZD.scala 39:21]
  assign _T_894 = _T_891[0]; // @[LZD.scala 39:30]
  assign _T_895 = ~ _T_894; // @[LZD.scala 39:27]
  assign _T_896 = _T_893 | _T_895; // @[LZD.scala 39:25]
  assign _T_897 = {_T_892,_T_896}; // @[Cat.scala 29:58]
  assign _T_898 = _T_890[1]; // @[Shift.scala 12:21]
  assign _T_899 = _T_897[1]; // @[Shift.scala 12:21]
  assign _T_900 = _T_898 | _T_899; // @[LZD.scala 49:16]
  assign _T_901 = ~ _T_899; // @[LZD.scala 49:27]
  assign _T_902 = _T_898 | _T_901; // @[LZD.scala 49:25]
  assign _T_903 = _T_890[0:0]; // @[LZD.scala 49:47]
  assign _T_904 = _T_897[0:0]; // @[LZD.scala 49:59]
  assign _T_905 = _T_898 ? _T_903 : _T_904; // @[LZD.scala 49:35]
  assign _T_907 = {_T_900,_T_902,_T_905}; // @[Cat.scala 29:58]
  assign _T_908 = _T_882[2]; // @[Shift.scala 12:21]
  assign _T_909 = _T_907[2]; // @[Shift.scala 12:21]
  assign _T_910 = _T_908 | _T_909; // @[LZD.scala 49:16]
  assign _T_911 = ~ _T_909; // @[LZD.scala 49:27]
  assign _T_912 = _T_908 | _T_911; // @[LZD.scala 49:25]
  assign _T_913 = _T_882[1:0]; // @[LZD.scala 49:47]
  assign _T_914 = _T_907[1:0]; // @[LZD.scala 49:59]
  assign _T_915 = _T_908 ? _T_913 : _T_914; // @[LZD.scala 49:35]
  assign _T_917 = {_T_910,_T_912,_T_915}; // @[Cat.scala 29:58]
  assign _T_918 = _T_856[7:0]; // @[LZD.scala 44:32]
  assign _T_919 = _T_918[7:4]; // @[LZD.scala 43:32]
  assign _T_920 = _T_919[3:2]; // @[LZD.scala 43:32]
  assign _T_921 = _T_920 != 2'h0; // @[LZD.scala 39:14]
  assign _T_922 = _T_920[1]; // @[LZD.scala 39:21]
  assign _T_923 = _T_920[0]; // @[LZD.scala 39:30]
  assign _T_924 = ~ _T_923; // @[LZD.scala 39:27]
  assign _T_925 = _T_922 | _T_924; // @[LZD.scala 39:25]
  assign _T_926 = {_T_921,_T_925}; // @[Cat.scala 29:58]
  assign _T_927 = _T_919[1:0]; // @[LZD.scala 44:32]
  assign _T_928 = _T_927 != 2'h0; // @[LZD.scala 39:14]
  assign _T_929 = _T_927[1]; // @[LZD.scala 39:21]
  assign _T_930 = _T_927[0]; // @[LZD.scala 39:30]
  assign _T_931 = ~ _T_930; // @[LZD.scala 39:27]
  assign _T_932 = _T_929 | _T_931; // @[LZD.scala 39:25]
  assign _T_933 = {_T_928,_T_932}; // @[Cat.scala 29:58]
  assign _T_934 = _T_926[1]; // @[Shift.scala 12:21]
  assign _T_935 = _T_933[1]; // @[Shift.scala 12:21]
  assign _T_936 = _T_934 | _T_935; // @[LZD.scala 49:16]
  assign _T_937 = ~ _T_935; // @[LZD.scala 49:27]
  assign _T_938 = _T_934 | _T_937; // @[LZD.scala 49:25]
  assign _T_939 = _T_926[0:0]; // @[LZD.scala 49:47]
  assign _T_940 = _T_933[0:0]; // @[LZD.scala 49:59]
  assign _T_941 = _T_934 ? _T_939 : _T_940; // @[LZD.scala 49:35]
  assign _T_943 = {_T_936,_T_938,_T_941}; // @[Cat.scala 29:58]
  assign _T_944 = _T_918[3:0]; // @[LZD.scala 44:32]
  assign _T_945 = _T_944[3:2]; // @[LZD.scala 43:32]
  assign _T_946 = _T_945 != 2'h0; // @[LZD.scala 39:14]
  assign _T_947 = _T_945[1]; // @[LZD.scala 39:21]
  assign _T_948 = _T_945[0]; // @[LZD.scala 39:30]
  assign _T_949 = ~ _T_948; // @[LZD.scala 39:27]
  assign _T_950 = _T_947 | _T_949; // @[LZD.scala 39:25]
  assign _T_951 = {_T_946,_T_950}; // @[Cat.scala 29:58]
  assign _T_952 = _T_944[1:0]; // @[LZD.scala 44:32]
  assign _T_953 = _T_952 != 2'h0; // @[LZD.scala 39:14]
  assign _T_954 = _T_952[1]; // @[LZD.scala 39:21]
  assign _T_955 = _T_952[0]; // @[LZD.scala 39:30]
  assign _T_956 = ~ _T_955; // @[LZD.scala 39:27]
  assign _T_957 = _T_954 | _T_956; // @[LZD.scala 39:25]
  assign _T_958 = {_T_953,_T_957}; // @[Cat.scala 29:58]
  assign _T_959 = _T_951[1]; // @[Shift.scala 12:21]
  assign _T_960 = _T_958[1]; // @[Shift.scala 12:21]
  assign _T_961 = _T_959 | _T_960; // @[LZD.scala 49:16]
  assign _T_962 = ~ _T_960; // @[LZD.scala 49:27]
  assign _T_963 = _T_959 | _T_962; // @[LZD.scala 49:25]
  assign _T_964 = _T_951[0:0]; // @[LZD.scala 49:47]
  assign _T_965 = _T_958[0:0]; // @[LZD.scala 49:59]
  assign _T_966 = _T_959 ? _T_964 : _T_965; // @[LZD.scala 49:35]
  assign _T_968 = {_T_961,_T_963,_T_966}; // @[Cat.scala 29:58]
  assign _T_969 = _T_943[2]; // @[Shift.scala 12:21]
  assign _T_970 = _T_968[2]; // @[Shift.scala 12:21]
  assign _T_971 = _T_969 | _T_970; // @[LZD.scala 49:16]
  assign _T_972 = ~ _T_970; // @[LZD.scala 49:27]
  assign _T_973 = _T_969 | _T_972; // @[LZD.scala 49:25]
  assign _T_974 = _T_943[1:0]; // @[LZD.scala 49:47]
  assign _T_975 = _T_968[1:0]; // @[LZD.scala 49:59]
  assign _T_976 = _T_969 ? _T_974 : _T_975; // @[LZD.scala 49:35]
  assign _T_978 = {_T_971,_T_973,_T_976}; // @[Cat.scala 29:58]
  assign _T_979 = _T_917[3]; // @[Shift.scala 12:21]
  assign _T_980 = _T_978[3]; // @[Shift.scala 12:21]
  assign _T_981 = _T_979 | _T_980; // @[LZD.scala 49:16]
  assign _T_982 = ~ _T_980; // @[LZD.scala 49:27]
  assign _T_983 = _T_979 | _T_982; // @[LZD.scala 49:25]
  assign _T_984 = _T_917[2:0]; // @[LZD.scala 49:47]
  assign _T_985 = _T_978[2:0]; // @[LZD.scala 49:59]
  assign _T_986 = _T_979 ? _T_984 : _T_985; // @[LZD.scala 49:35]
  assign _T_988 = {_T_981,_T_983,_T_986}; // @[Cat.scala 29:58]
  assign _T_989 = _T_855[15:0]; // @[LZD.scala 44:32]
  assign _T_990 = _T_989[15:8]; // @[LZD.scala 43:32]
  assign _T_991 = _T_990[7:4]; // @[LZD.scala 43:32]
  assign _T_992 = _T_991[3:2]; // @[LZD.scala 43:32]
  assign _T_993 = _T_992 != 2'h0; // @[LZD.scala 39:14]
  assign _T_994 = _T_992[1]; // @[LZD.scala 39:21]
  assign _T_995 = _T_992[0]; // @[LZD.scala 39:30]
  assign _T_996 = ~ _T_995; // @[LZD.scala 39:27]
  assign _T_997 = _T_994 | _T_996; // @[LZD.scala 39:25]
  assign _T_998 = {_T_993,_T_997}; // @[Cat.scala 29:58]
  assign _T_999 = _T_991[1:0]; // @[LZD.scala 44:32]
  assign _T_1000 = _T_999 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1001 = _T_999[1]; // @[LZD.scala 39:21]
  assign _T_1002 = _T_999[0]; // @[LZD.scala 39:30]
  assign _T_1003 = ~ _T_1002; // @[LZD.scala 39:27]
  assign _T_1004 = _T_1001 | _T_1003; // @[LZD.scala 39:25]
  assign _T_1005 = {_T_1000,_T_1004}; // @[Cat.scala 29:58]
  assign _T_1006 = _T_998[1]; // @[Shift.scala 12:21]
  assign _T_1007 = _T_1005[1]; // @[Shift.scala 12:21]
  assign _T_1008 = _T_1006 | _T_1007; // @[LZD.scala 49:16]
  assign _T_1009 = ~ _T_1007; // @[LZD.scala 49:27]
  assign _T_1010 = _T_1006 | _T_1009; // @[LZD.scala 49:25]
  assign _T_1011 = _T_998[0:0]; // @[LZD.scala 49:47]
  assign _T_1012 = _T_1005[0:0]; // @[LZD.scala 49:59]
  assign _T_1013 = _T_1006 ? _T_1011 : _T_1012; // @[LZD.scala 49:35]
  assign _T_1015 = {_T_1008,_T_1010,_T_1013}; // @[Cat.scala 29:58]
  assign _T_1016 = _T_990[3:0]; // @[LZD.scala 44:32]
  assign _T_1017 = _T_1016[3:2]; // @[LZD.scala 43:32]
  assign _T_1018 = _T_1017 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1019 = _T_1017[1]; // @[LZD.scala 39:21]
  assign _T_1020 = _T_1017[0]; // @[LZD.scala 39:30]
  assign _T_1021 = ~ _T_1020; // @[LZD.scala 39:27]
  assign _T_1022 = _T_1019 | _T_1021; // @[LZD.scala 39:25]
  assign _T_1023 = {_T_1018,_T_1022}; // @[Cat.scala 29:58]
  assign _T_1024 = _T_1016[1:0]; // @[LZD.scala 44:32]
  assign _T_1025 = _T_1024 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1026 = _T_1024[1]; // @[LZD.scala 39:21]
  assign _T_1027 = _T_1024[0]; // @[LZD.scala 39:30]
  assign _T_1028 = ~ _T_1027; // @[LZD.scala 39:27]
  assign _T_1029 = _T_1026 | _T_1028; // @[LZD.scala 39:25]
  assign _T_1030 = {_T_1025,_T_1029}; // @[Cat.scala 29:58]
  assign _T_1031 = _T_1023[1]; // @[Shift.scala 12:21]
  assign _T_1032 = _T_1030[1]; // @[Shift.scala 12:21]
  assign _T_1033 = _T_1031 | _T_1032; // @[LZD.scala 49:16]
  assign _T_1034 = ~ _T_1032; // @[LZD.scala 49:27]
  assign _T_1035 = _T_1031 | _T_1034; // @[LZD.scala 49:25]
  assign _T_1036 = _T_1023[0:0]; // @[LZD.scala 49:47]
  assign _T_1037 = _T_1030[0:0]; // @[LZD.scala 49:59]
  assign _T_1038 = _T_1031 ? _T_1036 : _T_1037; // @[LZD.scala 49:35]
  assign _T_1040 = {_T_1033,_T_1035,_T_1038}; // @[Cat.scala 29:58]
  assign _T_1041 = _T_1015[2]; // @[Shift.scala 12:21]
  assign _T_1042 = _T_1040[2]; // @[Shift.scala 12:21]
  assign _T_1043 = _T_1041 | _T_1042; // @[LZD.scala 49:16]
  assign _T_1044 = ~ _T_1042; // @[LZD.scala 49:27]
  assign _T_1045 = _T_1041 | _T_1044; // @[LZD.scala 49:25]
  assign _T_1046 = _T_1015[1:0]; // @[LZD.scala 49:47]
  assign _T_1047 = _T_1040[1:0]; // @[LZD.scala 49:59]
  assign _T_1048 = _T_1041 ? _T_1046 : _T_1047; // @[LZD.scala 49:35]
  assign _T_1050 = {_T_1043,_T_1045,_T_1048}; // @[Cat.scala 29:58]
  assign _T_1051 = _T_989[7:0]; // @[LZD.scala 44:32]
  assign _T_1052 = _T_1051[7:4]; // @[LZD.scala 43:32]
  assign _T_1053 = _T_1052[3:2]; // @[LZD.scala 43:32]
  assign _T_1054 = _T_1053 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1055 = _T_1053[1]; // @[LZD.scala 39:21]
  assign _T_1056 = _T_1053[0]; // @[LZD.scala 39:30]
  assign _T_1057 = ~ _T_1056; // @[LZD.scala 39:27]
  assign _T_1058 = _T_1055 | _T_1057; // @[LZD.scala 39:25]
  assign _T_1059 = {_T_1054,_T_1058}; // @[Cat.scala 29:58]
  assign _T_1060 = _T_1052[1:0]; // @[LZD.scala 44:32]
  assign _T_1061 = _T_1060 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1062 = _T_1060[1]; // @[LZD.scala 39:21]
  assign _T_1063 = _T_1060[0]; // @[LZD.scala 39:30]
  assign _T_1064 = ~ _T_1063; // @[LZD.scala 39:27]
  assign _T_1065 = _T_1062 | _T_1064; // @[LZD.scala 39:25]
  assign _T_1066 = {_T_1061,_T_1065}; // @[Cat.scala 29:58]
  assign _T_1067 = _T_1059[1]; // @[Shift.scala 12:21]
  assign _T_1068 = _T_1066[1]; // @[Shift.scala 12:21]
  assign _T_1069 = _T_1067 | _T_1068; // @[LZD.scala 49:16]
  assign _T_1070 = ~ _T_1068; // @[LZD.scala 49:27]
  assign _T_1071 = _T_1067 | _T_1070; // @[LZD.scala 49:25]
  assign _T_1072 = _T_1059[0:0]; // @[LZD.scala 49:47]
  assign _T_1073 = _T_1066[0:0]; // @[LZD.scala 49:59]
  assign _T_1074 = _T_1067 ? _T_1072 : _T_1073; // @[LZD.scala 49:35]
  assign _T_1076 = {_T_1069,_T_1071,_T_1074}; // @[Cat.scala 29:58]
  assign _T_1077 = _T_1051[3:0]; // @[LZD.scala 44:32]
  assign _T_1078 = _T_1077[3:2]; // @[LZD.scala 43:32]
  assign _T_1079 = _T_1078 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1080 = _T_1078[1]; // @[LZD.scala 39:21]
  assign _T_1081 = _T_1078[0]; // @[LZD.scala 39:30]
  assign _T_1082 = ~ _T_1081; // @[LZD.scala 39:27]
  assign _T_1083 = _T_1080 | _T_1082; // @[LZD.scala 39:25]
  assign _T_1084 = {_T_1079,_T_1083}; // @[Cat.scala 29:58]
  assign _T_1085 = _T_1077[1:0]; // @[LZD.scala 44:32]
  assign _T_1086 = _T_1085 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1087 = _T_1085[1]; // @[LZD.scala 39:21]
  assign _T_1088 = _T_1085[0]; // @[LZD.scala 39:30]
  assign _T_1089 = ~ _T_1088; // @[LZD.scala 39:27]
  assign _T_1090 = _T_1087 | _T_1089; // @[LZD.scala 39:25]
  assign _T_1091 = {_T_1086,_T_1090}; // @[Cat.scala 29:58]
  assign _T_1092 = _T_1084[1]; // @[Shift.scala 12:21]
  assign _T_1093 = _T_1091[1]; // @[Shift.scala 12:21]
  assign _T_1094 = _T_1092 | _T_1093; // @[LZD.scala 49:16]
  assign _T_1095 = ~ _T_1093; // @[LZD.scala 49:27]
  assign _T_1096 = _T_1092 | _T_1095; // @[LZD.scala 49:25]
  assign _T_1097 = _T_1084[0:0]; // @[LZD.scala 49:47]
  assign _T_1098 = _T_1091[0:0]; // @[LZD.scala 49:59]
  assign _T_1099 = _T_1092 ? _T_1097 : _T_1098; // @[LZD.scala 49:35]
  assign _T_1101 = {_T_1094,_T_1096,_T_1099}; // @[Cat.scala 29:58]
  assign _T_1102 = _T_1076[2]; // @[Shift.scala 12:21]
  assign _T_1103 = _T_1101[2]; // @[Shift.scala 12:21]
  assign _T_1104 = _T_1102 | _T_1103; // @[LZD.scala 49:16]
  assign _T_1105 = ~ _T_1103; // @[LZD.scala 49:27]
  assign _T_1106 = _T_1102 | _T_1105; // @[LZD.scala 49:25]
  assign _T_1107 = _T_1076[1:0]; // @[LZD.scala 49:47]
  assign _T_1108 = _T_1101[1:0]; // @[LZD.scala 49:59]
  assign _T_1109 = _T_1102 ? _T_1107 : _T_1108; // @[LZD.scala 49:35]
  assign _T_1111 = {_T_1104,_T_1106,_T_1109}; // @[Cat.scala 29:58]
  assign _T_1112 = _T_1050[3]; // @[Shift.scala 12:21]
  assign _T_1113 = _T_1111[3]; // @[Shift.scala 12:21]
  assign _T_1114 = _T_1112 | _T_1113; // @[LZD.scala 49:16]
  assign _T_1115 = ~ _T_1113; // @[LZD.scala 49:27]
  assign _T_1116 = _T_1112 | _T_1115; // @[LZD.scala 49:25]
  assign _T_1117 = _T_1050[2:0]; // @[LZD.scala 49:47]
  assign _T_1118 = _T_1111[2:0]; // @[LZD.scala 49:59]
  assign _T_1119 = _T_1112 ? _T_1117 : _T_1118; // @[LZD.scala 49:35]
  assign _T_1121 = {_T_1114,_T_1116,_T_1119}; // @[Cat.scala 29:58]
  assign _T_1122 = _T_988[4]; // @[Shift.scala 12:21]
  assign _T_1123 = _T_1121[4]; // @[Shift.scala 12:21]
  assign _T_1124 = _T_1122 | _T_1123; // @[LZD.scala 49:16]
  assign _T_1125 = ~ _T_1123; // @[LZD.scala 49:27]
  assign _T_1126 = _T_1122 | _T_1125; // @[LZD.scala 49:25]
  assign _T_1127 = _T_988[3:0]; // @[LZD.scala 49:47]
  assign _T_1128 = _T_1121[3:0]; // @[LZD.scala 49:59]
  assign _T_1129 = _T_1122 ? _T_1127 : _T_1128; // @[LZD.scala 49:35]
  assign _T_1131 = {_T_1124,_T_1126,_T_1129}; // @[Cat.scala 29:58]
  assign _T_1132 = _T_854[5]; // @[Shift.scala 12:21]
  assign _T_1133 = _T_1131[5]; // @[Shift.scala 12:21]
  assign _T_1134 = _T_1132 | _T_1133; // @[LZD.scala 49:16]
  assign _T_1135 = ~ _T_1133; // @[LZD.scala 49:27]
  assign _T_1136 = _T_1132 | _T_1135; // @[LZD.scala 49:25]
  assign _T_1137 = _T_854[4:0]; // @[LZD.scala 49:47]
  assign _T_1138 = _T_1131[4:0]; // @[LZD.scala 49:59]
  assign _T_1139 = _T_1132 ? _T_1137 : _T_1138; // @[LZD.scala 49:35]
  assign _T_1141 = {_T_1134,_T_1136,_T_1139}; // @[Cat.scala 29:58]
  assign _T_1142 = _T_576[6]; // @[Shift.scala 12:21]
  assign _T_1143 = _T_1141[6]; // @[Shift.scala 12:21]
  assign _T_1144 = _T_1142 | _T_1143; // @[LZD.scala 49:16]
  assign _T_1145 = ~ _T_1143; // @[LZD.scala 49:27]
  assign _T_1146 = _T_1142 | _T_1145; // @[LZD.scala 49:25]
  assign _T_1147 = _T_576[5:0]; // @[LZD.scala 49:47]
  assign _T_1148 = _T_1141[5:0]; // @[LZD.scala 49:59]
  assign _T_1149 = _T_1142 ? _T_1147 : _T_1148; // @[LZD.scala 49:35]
  assign _T_1151 = {_T_1144,_T_1146,_T_1149}; // @[Cat.scala 29:58]
  assign _T_1152 = _T_10[127:0]; // @[LZD.scala 44:32]
  assign _T_1153 = _T_1152[127:64]; // @[LZD.scala 43:32]
  assign _T_1154 = _T_1153[63:32]; // @[LZD.scala 43:32]
  assign _T_1155 = _T_1154[31:16]; // @[LZD.scala 43:32]
  assign _T_1156 = _T_1155[15:8]; // @[LZD.scala 43:32]
  assign _T_1157 = _T_1156[7:4]; // @[LZD.scala 43:32]
  assign _T_1158 = _T_1157[3:2]; // @[LZD.scala 43:32]
  assign _T_1159 = _T_1158 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1160 = _T_1158[1]; // @[LZD.scala 39:21]
  assign _T_1161 = _T_1158[0]; // @[LZD.scala 39:30]
  assign _T_1162 = ~ _T_1161; // @[LZD.scala 39:27]
  assign _T_1163 = _T_1160 | _T_1162; // @[LZD.scala 39:25]
  assign _T_1164 = {_T_1159,_T_1163}; // @[Cat.scala 29:58]
  assign _T_1165 = _T_1157[1:0]; // @[LZD.scala 44:32]
  assign _T_1166 = _T_1165 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1167 = _T_1165[1]; // @[LZD.scala 39:21]
  assign _T_1168 = _T_1165[0]; // @[LZD.scala 39:30]
  assign _T_1169 = ~ _T_1168; // @[LZD.scala 39:27]
  assign _T_1170 = _T_1167 | _T_1169; // @[LZD.scala 39:25]
  assign _T_1171 = {_T_1166,_T_1170}; // @[Cat.scala 29:58]
  assign _T_1172 = _T_1164[1]; // @[Shift.scala 12:21]
  assign _T_1173 = _T_1171[1]; // @[Shift.scala 12:21]
  assign _T_1174 = _T_1172 | _T_1173; // @[LZD.scala 49:16]
  assign _T_1175 = ~ _T_1173; // @[LZD.scala 49:27]
  assign _T_1176 = _T_1172 | _T_1175; // @[LZD.scala 49:25]
  assign _T_1177 = _T_1164[0:0]; // @[LZD.scala 49:47]
  assign _T_1178 = _T_1171[0:0]; // @[LZD.scala 49:59]
  assign _T_1179 = _T_1172 ? _T_1177 : _T_1178; // @[LZD.scala 49:35]
  assign _T_1181 = {_T_1174,_T_1176,_T_1179}; // @[Cat.scala 29:58]
  assign _T_1182 = _T_1156[3:0]; // @[LZD.scala 44:32]
  assign _T_1183 = _T_1182[3:2]; // @[LZD.scala 43:32]
  assign _T_1184 = _T_1183 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1185 = _T_1183[1]; // @[LZD.scala 39:21]
  assign _T_1186 = _T_1183[0]; // @[LZD.scala 39:30]
  assign _T_1187 = ~ _T_1186; // @[LZD.scala 39:27]
  assign _T_1188 = _T_1185 | _T_1187; // @[LZD.scala 39:25]
  assign _T_1189 = {_T_1184,_T_1188}; // @[Cat.scala 29:58]
  assign _T_1190 = _T_1182[1:0]; // @[LZD.scala 44:32]
  assign _T_1191 = _T_1190 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1192 = _T_1190[1]; // @[LZD.scala 39:21]
  assign _T_1193 = _T_1190[0]; // @[LZD.scala 39:30]
  assign _T_1194 = ~ _T_1193; // @[LZD.scala 39:27]
  assign _T_1195 = _T_1192 | _T_1194; // @[LZD.scala 39:25]
  assign _T_1196 = {_T_1191,_T_1195}; // @[Cat.scala 29:58]
  assign _T_1197 = _T_1189[1]; // @[Shift.scala 12:21]
  assign _T_1198 = _T_1196[1]; // @[Shift.scala 12:21]
  assign _T_1199 = _T_1197 | _T_1198; // @[LZD.scala 49:16]
  assign _T_1200 = ~ _T_1198; // @[LZD.scala 49:27]
  assign _T_1201 = _T_1197 | _T_1200; // @[LZD.scala 49:25]
  assign _T_1202 = _T_1189[0:0]; // @[LZD.scala 49:47]
  assign _T_1203 = _T_1196[0:0]; // @[LZD.scala 49:59]
  assign _T_1204 = _T_1197 ? _T_1202 : _T_1203; // @[LZD.scala 49:35]
  assign _T_1206 = {_T_1199,_T_1201,_T_1204}; // @[Cat.scala 29:58]
  assign _T_1207 = _T_1181[2]; // @[Shift.scala 12:21]
  assign _T_1208 = _T_1206[2]; // @[Shift.scala 12:21]
  assign _T_1209 = _T_1207 | _T_1208; // @[LZD.scala 49:16]
  assign _T_1210 = ~ _T_1208; // @[LZD.scala 49:27]
  assign _T_1211 = _T_1207 | _T_1210; // @[LZD.scala 49:25]
  assign _T_1212 = _T_1181[1:0]; // @[LZD.scala 49:47]
  assign _T_1213 = _T_1206[1:0]; // @[LZD.scala 49:59]
  assign _T_1214 = _T_1207 ? _T_1212 : _T_1213; // @[LZD.scala 49:35]
  assign _T_1216 = {_T_1209,_T_1211,_T_1214}; // @[Cat.scala 29:58]
  assign _T_1217 = _T_1155[7:0]; // @[LZD.scala 44:32]
  assign _T_1218 = _T_1217[7:4]; // @[LZD.scala 43:32]
  assign _T_1219 = _T_1218[3:2]; // @[LZD.scala 43:32]
  assign _T_1220 = _T_1219 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1221 = _T_1219[1]; // @[LZD.scala 39:21]
  assign _T_1222 = _T_1219[0]; // @[LZD.scala 39:30]
  assign _T_1223 = ~ _T_1222; // @[LZD.scala 39:27]
  assign _T_1224 = _T_1221 | _T_1223; // @[LZD.scala 39:25]
  assign _T_1225 = {_T_1220,_T_1224}; // @[Cat.scala 29:58]
  assign _T_1226 = _T_1218[1:0]; // @[LZD.scala 44:32]
  assign _T_1227 = _T_1226 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1228 = _T_1226[1]; // @[LZD.scala 39:21]
  assign _T_1229 = _T_1226[0]; // @[LZD.scala 39:30]
  assign _T_1230 = ~ _T_1229; // @[LZD.scala 39:27]
  assign _T_1231 = _T_1228 | _T_1230; // @[LZD.scala 39:25]
  assign _T_1232 = {_T_1227,_T_1231}; // @[Cat.scala 29:58]
  assign _T_1233 = _T_1225[1]; // @[Shift.scala 12:21]
  assign _T_1234 = _T_1232[1]; // @[Shift.scala 12:21]
  assign _T_1235 = _T_1233 | _T_1234; // @[LZD.scala 49:16]
  assign _T_1236 = ~ _T_1234; // @[LZD.scala 49:27]
  assign _T_1237 = _T_1233 | _T_1236; // @[LZD.scala 49:25]
  assign _T_1238 = _T_1225[0:0]; // @[LZD.scala 49:47]
  assign _T_1239 = _T_1232[0:0]; // @[LZD.scala 49:59]
  assign _T_1240 = _T_1233 ? _T_1238 : _T_1239; // @[LZD.scala 49:35]
  assign _T_1242 = {_T_1235,_T_1237,_T_1240}; // @[Cat.scala 29:58]
  assign _T_1243 = _T_1217[3:0]; // @[LZD.scala 44:32]
  assign _T_1244 = _T_1243[3:2]; // @[LZD.scala 43:32]
  assign _T_1245 = _T_1244 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1246 = _T_1244[1]; // @[LZD.scala 39:21]
  assign _T_1247 = _T_1244[0]; // @[LZD.scala 39:30]
  assign _T_1248 = ~ _T_1247; // @[LZD.scala 39:27]
  assign _T_1249 = _T_1246 | _T_1248; // @[LZD.scala 39:25]
  assign _T_1250 = {_T_1245,_T_1249}; // @[Cat.scala 29:58]
  assign _T_1251 = _T_1243[1:0]; // @[LZD.scala 44:32]
  assign _T_1252 = _T_1251 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1253 = _T_1251[1]; // @[LZD.scala 39:21]
  assign _T_1254 = _T_1251[0]; // @[LZD.scala 39:30]
  assign _T_1255 = ~ _T_1254; // @[LZD.scala 39:27]
  assign _T_1256 = _T_1253 | _T_1255; // @[LZD.scala 39:25]
  assign _T_1257 = {_T_1252,_T_1256}; // @[Cat.scala 29:58]
  assign _T_1258 = _T_1250[1]; // @[Shift.scala 12:21]
  assign _T_1259 = _T_1257[1]; // @[Shift.scala 12:21]
  assign _T_1260 = _T_1258 | _T_1259; // @[LZD.scala 49:16]
  assign _T_1261 = ~ _T_1259; // @[LZD.scala 49:27]
  assign _T_1262 = _T_1258 | _T_1261; // @[LZD.scala 49:25]
  assign _T_1263 = _T_1250[0:0]; // @[LZD.scala 49:47]
  assign _T_1264 = _T_1257[0:0]; // @[LZD.scala 49:59]
  assign _T_1265 = _T_1258 ? _T_1263 : _T_1264; // @[LZD.scala 49:35]
  assign _T_1267 = {_T_1260,_T_1262,_T_1265}; // @[Cat.scala 29:58]
  assign _T_1268 = _T_1242[2]; // @[Shift.scala 12:21]
  assign _T_1269 = _T_1267[2]; // @[Shift.scala 12:21]
  assign _T_1270 = _T_1268 | _T_1269; // @[LZD.scala 49:16]
  assign _T_1271 = ~ _T_1269; // @[LZD.scala 49:27]
  assign _T_1272 = _T_1268 | _T_1271; // @[LZD.scala 49:25]
  assign _T_1273 = _T_1242[1:0]; // @[LZD.scala 49:47]
  assign _T_1274 = _T_1267[1:0]; // @[LZD.scala 49:59]
  assign _T_1275 = _T_1268 ? _T_1273 : _T_1274; // @[LZD.scala 49:35]
  assign _T_1277 = {_T_1270,_T_1272,_T_1275}; // @[Cat.scala 29:58]
  assign _T_1278 = _T_1216[3]; // @[Shift.scala 12:21]
  assign _T_1279 = _T_1277[3]; // @[Shift.scala 12:21]
  assign _T_1280 = _T_1278 | _T_1279; // @[LZD.scala 49:16]
  assign _T_1281 = ~ _T_1279; // @[LZD.scala 49:27]
  assign _T_1282 = _T_1278 | _T_1281; // @[LZD.scala 49:25]
  assign _T_1283 = _T_1216[2:0]; // @[LZD.scala 49:47]
  assign _T_1284 = _T_1277[2:0]; // @[LZD.scala 49:59]
  assign _T_1285 = _T_1278 ? _T_1283 : _T_1284; // @[LZD.scala 49:35]
  assign _T_1287 = {_T_1280,_T_1282,_T_1285}; // @[Cat.scala 29:58]
  assign _T_1288 = _T_1154[15:0]; // @[LZD.scala 44:32]
  assign _T_1289 = _T_1288[15:8]; // @[LZD.scala 43:32]
  assign _T_1290 = _T_1289[7:4]; // @[LZD.scala 43:32]
  assign _T_1291 = _T_1290[3:2]; // @[LZD.scala 43:32]
  assign _T_1292 = _T_1291 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1293 = _T_1291[1]; // @[LZD.scala 39:21]
  assign _T_1294 = _T_1291[0]; // @[LZD.scala 39:30]
  assign _T_1295 = ~ _T_1294; // @[LZD.scala 39:27]
  assign _T_1296 = _T_1293 | _T_1295; // @[LZD.scala 39:25]
  assign _T_1297 = {_T_1292,_T_1296}; // @[Cat.scala 29:58]
  assign _T_1298 = _T_1290[1:0]; // @[LZD.scala 44:32]
  assign _T_1299 = _T_1298 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1300 = _T_1298[1]; // @[LZD.scala 39:21]
  assign _T_1301 = _T_1298[0]; // @[LZD.scala 39:30]
  assign _T_1302 = ~ _T_1301; // @[LZD.scala 39:27]
  assign _T_1303 = _T_1300 | _T_1302; // @[LZD.scala 39:25]
  assign _T_1304 = {_T_1299,_T_1303}; // @[Cat.scala 29:58]
  assign _T_1305 = _T_1297[1]; // @[Shift.scala 12:21]
  assign _T_1306 = _T_1304[1]; // @[Shift.scala 12:21]
  assign _T_1307 = _T_1305 | _T_1306; // @[LZD.scala 49:16]
  assign _T_1308 = ~ _T_1306; // @[LZD.scala 49:27]
  assign _T_1309 = _T_1305 | _T_1308; // @[LZD.scala 49:25]
  assign _T_1310 = _T_1297[0:0]; // @[LZD.scala 49:47]
  assign _T_1311 = _T_1304[0:0]; // @[LZD.scala 49:59]
  assign _T_1312 = _T_1305 ? _T_1310 : _T_1311; // @[LZD.scala 49:35]
  assign _T_1314 = {_T_1307,_T_1309,_T_1312}; // @[Cat.scala 29:58]
  assign _T_1315 = _T_1289[3:0]; // @[LZD.scala 44:32]
  assign _T_1316 = _T_1315[3:2]; // @[LZD.scala 43:32]
  assign _T_1317 = _T_1316 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1318 = _T_1316[1]; // @[LZD.scala 39:21]
  assign _T_1319 = _T_1316[0]; // @[LZD.scala 39:30]
  assign _T_1320 = ~ _T_1319; // @[LZD.scala 39:27]
  assign _T_1321 = _T_1318 | _T_1320; // @[LZD.scala 39:25]
  assign _T_1322 = {_T_1317,_T_1321}; // @[Cat.scala 29:58]
  assign _T_1323 = _T_1315[1:0]; // @[LZD.scala 44:32]
  assign _T_1324 = _T_1323 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1325 = _T_1323[1]; // @[LZD.scala 39:21]
  assign _T_1326 = _T_1323[0]; // @[LZD.scala 39:30]
  assign _T_1327 = ~ _T_1326; // @[LZD.scala 39:27]
  assign _T_1328 = _T_1325 | _T_1327; // @[LZD.scala 39:25]
  assign _T_1329 = {_T_1324,_T_1328}; // @[Cat.scala 29:58]
  assign _T_1330 = _T_1322[1]; // @[Shift.scala 12:21]
  assign _T_1331 = _T_1329[1]; // @[Shift.scala 12:21]
  assign _T_1332 = _T_1330 | _T_1331; // @[LZD.scala 49:16]
  assign _T_1333 = ~ _T_1331; // @[LZD.scala 49:27]
  assign _T_1334 = _T_1330 | _T_1333; // @[LZD.scala 49:25]
  assign _T_1335 = _T_1322[0:0]; // @[LZD.scala 49:47]
  assign _T_1336 = _T_1329[0:0]; // @[LZD.scala 49:59]
  assign _T_1337 = _T_1330 ? _T_1335 : _T_1336; // @[LZD.scala 49:35]
  assign _T_1339 = {_T_1332,_T_1334,_T_1337}; // @[Cat.scala 29:58]
  assign _T_1340 = _T_1314[2]; // @[Shift.scala 12:21]
  assign _T_1341 = _T_1339[2]; // @[Shift.scala 12:21]
  assign _T_1342 = _T_1340 | _T_1341; // @[LZD.scala 49:16]
  assign _T_1343 = ~ _T_1341; // @[LZD.scala 49:27]
  assign _T_1344 = _T_1340 | _T_1343; // @[LZD.scala 49:25]
  assign _T_1345 = _T_1314[1:0]; // @[LZD.scala 49:47]
  assign _T_1346 = _T_1339[1:0]; // @[LZD.scala 49:59]
  assign _T_1347 = _T_1340 ? _T_1345 : _T_1346; // @[LZD.scala 49:35]
  assign _T_1349 = {_T_1342,_T_1344,_T_1347}; // @[Cat.scala 29:58]
  assign _T_1350 = _T_1288[7:0]; // @[LZD.scala 44:32]
  assign _T_1351 = _T_1350[7:4]; // @[LZD.scala 43:32]
  assign _T_1352 = _T_1351[3:2]; // @[LZD.scala 43:32]
  assign _T_1353 = _T_1352 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1354 = _T_1352[1]; // @[LZD.scala 39:21]
  assign _T_1355 = _T_1352[0]; // @[LZD.scala 39:30]
  assign _T_1356 = ~ _T_1355; // @[LZD.scala 39:27]
  assign _T_1357 = _T_1354 | _T_1356; // @[LZD.scala 39:25]
  assign _T_1358 = {_T_1353,_T_1357}; // @[Cat.scala 29:58]
  assign _T_1359 = _T_1351[1:0]; // @[LZD.scala 44:32]
  assign _T_1360 = _T_1359 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1361 = _T_1359[1]; // @[LZD.scala 39:21]
  assign _T_1362 = _T_1359[0]; // @[LZD.scala 39:30]
  assign _T_1363 = ~ _T_1362; // @[LZD.scala 39:27]
  assign _T_1364 = _T_1361 | _T_1363; // @[LZD.scala 39:25]
  assign _T_1365 = {_T_1360,_T_1364}; // @[Cat.scala 29:58]
  assign _T_1366 = _T_1358[1]; // @[Shift.scala 12:21]
  assign _T_1367 = _T_1365[1]; // @[Shift.scala 12:21]
  assign _T_1368 = _T_1366 | _T_1367; // @[LZD.scala 49:16]
  assign _T_1369 = ~ _T_1367; // @[LZD.scala 49:27]
  assign _T_1370 = _T_1366 | _T_1369; // @[LZD.scala 49:25]
  assign _T_1371 = _T_1358[0:0]; // @[LZD.scala 49:47]
  assign _T_1372 = _T_1365[0:0]; // @[LZD.scala 49:59]
  assign _T_1373 = _T_1366 ? _T_1371 : _T_1372; // @[LZD.scala 49:35]
  assign _T_1375 = {_T_1368,_T_1370,_T_1373}; // @[Cat.scala 29:58]
  assign _T_1376 = _T_1350[3:0]; // @[LZD.scala 44:32]
  assign _T_1377 = _T_1376[3:2]; // @[LZD.scala 43:32]
  assign _T_1378 = _T_1377 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1379 = _T_1377[1]; // @[LZD.scala 39:21]
  assign _T_1380 = _T_1377[0]; // @[LZD.scala 39:30]
  assign _T_1381 = ~ _T_1380; // @[LZD.scala 39:27]
  assign _T_1382 = _T_1379 | _T_1381; // @[LZD.scala 39:25]
  assign _T_1383 = {_T_1378,_T_1382}; // @[Cat.scala 29:58]
  assign _T_1384 = _T_1376[1:0]; // @[LZD.scala 44:32]
  assign _T_1385 = _T_1384 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1386 = _T_1384[1]; // @[LZD.scala 39:21]
  assign _T_1387 = _T_1384[0]; // @[LZD.scala 39:30]
  assign _T_1388 = ~ _T_1387; // @[LZD.scala 39:27]
  assign _T_1389 = _T_1386 | _T_1388; // @[LZD.scala 39:25]
  assign _T_1390 = {_T_1385,_T_1389}; // @[Cat.scala 29:58]
  assign _T_1391 = _T_1383[1]; // @[Shift.scala 12:21]
  assign _T_1392 = _T_1390[1]; // @[Shift.scala 12:21]
  assign _T_1393 = _T_1391 | _T_1392; // @[LZD.scala 49:16]
  assign _T_1394 = ~ _T_1392; // @[LZD.scala 49:27]
  assign _T_1395 = _T_1391 | _T_1394; // @[LZD.scala 49:25]
  assign _T_1396 = _T_1383[0:0]; // @[LZD.scala 49:47]
  assign _T_1397 = _T_1390[0:0]; // @[LZD.scala 49:59]
  assign _T_1398 = _T_1391 ? _T_1396 : _T_1397; // @[LZD.scala 49:35]
  assign _T_1400 = {_T_1393,_T_1395,_T_1398}; // @[Cat.scala 29:58]
  assign _T_1401 = _T_1375[2]; // @[Shift.scala 12:21]
  assign _T_1402 = _T_1400[2]; // @[Shift.scala 12:21]
  assign _T_1403 = _T_1401 | _T_1402; // @[LZD.scala 49:16]
  assign _T_1404 = ~ _T_1402; // @[LZD.scala 49:27]
  assign _T_1405 = _T_1401 | _T_1404; // @[LZD.scala 49:25]
  assign _T_1406 = _T_1375[1:0]; // @[LZD.scala 49:47]
  assign _T_1407 = _T_1400[1:0]; // @[LZD.scala 49:59]
  assign _T_1408 = _T_1401 ? _T_1406 : _T_1407; // @[LZD.scala 49:35]
  assign _T_1410 = {_T_1403,_T_1405,_T_1408}; // @[Cat.scala 29:58]
  assign _T_1411 = _T_1349[3]; // @[Shift.scala 12:21]
  assign _T_1412 = _T_1410[3]; // @[Shift.scala 12:21]
  assign _T_1413 = _T_1411 | _T_1412; // @[LZD.scala 49:16]
  assign _T_1414 = ~ _T_1412; // @[LZD.scala 49:27]
  assign _T_1415 = _T_1411 | _T_1414; // @[LZD.scala 49:25]
  assign _T_1416 = _T_1349[2:0]; // @[LZD.scala 49:47]
  assign _T_1417 = _T_1410[2:0]; // @[LZD.scala 49:59]
  assign _T_1418 = _T_1411 ? _T_1416 : _T_1417; // @[LZD.scala 49:35]
  assign _T_1420 = {_T_1413,_T_1415,_T_1418}; // @[Cat.scala 29:58]
  assign _T_1421 = _T_1287[4]; // @[Shift.scala 12:21]
  assign _T_1422 = _T_1420[4]; // @[Shift.scala 12:21]
  assign _T_1423 = _T_1421 | _T_1422; // @[LZD.scala 49:16]
  assign _T_1424 = ~ _T_1422; // @[LZD.scala 49:27]
  assign _T_1425 = _T_1421 | _T_1424; // @[LZD.scala 49:25]
  assign _T_1426 = _T_1287[3:0]; // @[LZD.scala 49:47]
  assign _T_1427 = _T_1420[3:0]; // @[LZD.scala 49:59]
  assign _T_1428 = _T_1421 ? _T_1426 : _T_1427; // @[LZD.scala 49:35]
  assign _T_1430 = {_T_1423,_T_1425,_T_1428}; // @[Cat.scala 29:58]
  assign _T_1431 = _T_1153[31:0]; // @[LZD.scala 44:32]
  assign _T_1432 = _T_1431[31:16]; // @[LZD.scala 43:32]
  assign _T_1433 = _T_1432[15:8]; // @[LZD.scala 43:32]
  assign _T_1434 = _T_1433[7:4]; // @[LZD.scala 43:32]
  assign _T_1435 = _T_1434[3:2]; // @[LZD.scala 43:32]
  assign _T_1436 = _T_1435 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1437 = _T_1435[1]; // @[LZD.scala 39:21]
  assign _T_1438 = _T_1435[0]; // @[LZD.scala 39:30]
  assign _T_1439 = ~ _T_1438; // @[LZD.scala 39:27]
  assign _T_1440 = _T_1437 | _T_1439; // @[LZD.scala 39:25]
  assign _T_1441 = {_T_1436,_T_1440}; // @[Cat.scala 29:58]
  assign _T_1442 = _T_1434[1:0]; // @[LZD.scala 44:32]
  assign _T_1443 = _T_1442 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1444 = _T_1442[1]; // @[LZD.scala 39:21]
  assign _T_1445 = _T_1442[0]; // @[LZD.scala 39:30]
  assign _T_1446 = ~ _T_1445; // @[LZD.scala 39:27]
  assign _T_1447 = _T_1444 | _T_1446; // @[LZD.scala 39:25]
  assign _T_1448 = {_T_1443,_T_1447}; // @[Cat.scala 29:58]
  assign _T_1449 = _T_1441[1]; // @[Shift.scala 12:21]
  assign _T_1450 = _T_1448[1]; // @[Shift.scala 12:21]
  assign _T_1451 = _T_1449 | _T_1450; // @[LZD.scala 49:16]
  assign _T_1452 = ~ _T_1450; // @[LZD.scala 49:27]
  assign _T_1453 = _T_1449 | _T_1452; // @[LZD.scala 49:25]
  assign _T_1454 = _T_1441[0:0]; // @[LZD.scala 49:47]
  assign _T_1455 = _T_1448[0:0]; // @[LZD.scala 49:59]
  assign _T_1456 = _T_1449 ? _T_1454 : _T_1455; // @[LZD.scala 49:35]
  assign _T_1458 = {_T_1451,_T_1453,_T_1456}; // @[Cat.scala 29:58]
  assign _T_1459 = _T_1433[3:0]; // @[LZD.scala 44:32]
  assign _T_1460 = _T_1459[3:2]; // @[LZD.scala 43:32]
  assign _T_1461 = _T_1460 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1462 = _T_1460[1]; // @[LZD.scala 39:21]
  assign _T_1463 = _T_1460[0]; // @[LZD.scala 39:30]
  assign _T_1464 = ~ _T_1463; // @[LZD.scala 39:27]
  assign _T_1465 = _T_1462 | _T_1464; // @[LZD.scala 39:25]
  assign _T_1466 = {_T_1461,_T_1465}; // @[Cat.scala 29:58]
  assign _T_1467 = _T_1459[1:0]; // @[LZD.scala 44:32]
  assign _T_1468 = _T_1467 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1469 = _T_1467[1]; // @[LZD.scala 39:21]
  assign _T_1470 = _T_1467[0]; // @[LZD.scala 39:30]
  assign _T_1471 = ~ _T_1470; // @[LZD.scala 39:27]
  assign _T_1472 = _T_1469 | _T_1471; // @[LZD.scala 39:25]
  assign _T_1473 = {_T_1468,_T_1472}; // @[Cat.scala 29:58]
  assign _T_1474 = _T_1466[1]; // @[Shift.scala 12:21]
  assign _T_1475 = _T_1473[1]; // @[Shift.scala 12:21]
  assign _T_1476 = _T_1474 | _T_1475; // @[LZD.scala 49:16]
  assign _T_1477 = ~ _T_1475; // @[LZD.scala 49:27]
  assign _T_1478 = _T_1474 | _T_1477; // @[LZD.scala 49:25]
  assign _T_1479 = _T_1466[0:0]; // @[LZD.scala 49:47]
  assign _T_1480 = _T_1473[0:0]; // @[LZD.scala 49:59]
  assign _T_1481 = _T_1474 ? _T_1479 : _T_1480; // @[LZD.scala 49:35]
  assign _T_1483 = {_T_1476,_T_1478,_T_1481}; // @[Cat.scala 29:58]
  assign _T_1484 = _T_1458[2]; // @[Shift.scala 12:21]
  assign _T_1485 = _T_1483[2]; // @[Shift.scala 12:21]
  assign _T_1486 = _T_1484 | _T_1485; // @[LZD.scala 49:16]
  assign _T_1487 = ~ _T_1485; // @[LZD.scala 49:27]
  assign _T_1488 = _T_1484 | _T_1487; // @[LZD.scala 49:25]
  assign _T_1489 = _T_1458[1:0]; // @[LZD.scala 49:47]
  assign _T_1490 = _T_1483[1:0]; // @[LZD.scala 49:59]
  assign _T_1491 = _T_1484 ? _T_1489 : _T_1490; // @[LZD.scala 49:35]
  assign _T_1493 = {_T_1486,_T_1488,_T_1491}; // @[Cat.scala 29:58]
  assign _T_1494 = _T_1432[7:0]; // @[LZD.scala 44:32]
  assign _T_1495 = _T_1494[7:4]; // @[LZD.scala 43:32]
  assign _T_1496 = _T_1495[3:2]; // @[LZD.scala 43:32]
  assign _T_1497 = _T_1496 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1498 = _T_1496[1]; // @[LZD.scala 39:21]
  assign _T_1499 = _T_1496[0]; // @[LZD.scala 39:30]
  assign _T_1500 = ~ _T_1499; // @[LZD.scala 39:27]
  assign _T_1501 = _T_1498 | _T_1500; // @[LZD.scala 39:25]
  assign _T_1502 = {_T_1497,_T_1501}; // @[Cat.scala 29:58]
  assign _T_1503 = _T_1495[1:0]; // @[LZD.scala 44:32]
  assign _T_1504 = _T_1503 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1505 = _T_1503[1]; // @[LZD.scala 39:21]
  assign _T_1506 = _T_1503[0]; // @[LZD.scala 39:30]
  assign _T_1507 = ~ _T_1506; // @[LZD.scala 39:27]
  assign _T_1508 = _T_1505 | _T_1507; // @[LZD.scala 39:25]
  assign _T_1509 = {_T_1504,_T_1508}; // @[Cat.scala 29:58]
  assign _T_1510 = _T_1502[1]; // @[Shift.scala 12:21]
  assign _T_1511 = _T_1509[1]; // @[Shift.scala 12:21]
  assign _T_1512 = _T_1510 | _T_1511; // @[LZD.scala 49:16]
  assign _T_1513 = ~ _T_1511; // @[LZD.scala 49:27]
  assign _T_1514 = _T_1510 | _T_1513; // @[LZD.scala 49:25]
  assign _T_1515 = _T_1502[0:0]; // @[LZD.scala 49:47]
  assign _T_1516 = _T_1509[0:0]; // @[LZD.scala 49:59]
  assign _T_1517 = _T_1510 ? _T_1515 : _T_1516; // @[LZD.scala 49:35]
  assign _T_1519 = {_T_1512,_T_1514,_T_1517}; // @[Cat.scala 29:58]
  assign _T_1520 = _T_1494[3:0]; // @[LZD.scala 44:32]
  assign _T_1521 = _T_1520[3:2]; // @[LZD.scala 43:32]
  assign _T_1522 = _T_1521 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1523 = _T_1521[1]; // @[LZD.scala 39:21]
  assign _T_1524 = _T_1521[0]; // @[LZD.scala 39:30]
  assign _T_1525 = ~ _T_1524; // @[LZD.scala 39:27]
  assign _T_1526 = _T_1523 | _T_1525; // @[LZD.scala 39:25]
  assign _T_1527 = {_T_1522,_T_1526}; // @[Cat.scala 29:58]
  assign _T_1528 = _T_1520[1:0]; // @[LZD.scala 44:32]
  assign _T_1529 = _T_1528 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1530 = _T_1528[1]; // @[LZD.scala 39:21]
  assign _T_1531 = _T_1528[0]; // @[LZD.scala 39:30]
  assign _T_1532 = ~ _T_1531; // @[LZD.scala 39:27]
  assign _T_1533 = _T_1530 | _T_1532; // @[LZD.scala 39:25]
  assign _T_1534 = {_T_1529,_T_1533}; // @[Cat.scala 29:58]
  assign _T_1535 = _T_1527[1]; // @[Shift.scala 12:21]
  assign _T_1536 = _T_1534[1]; // @[Shift.scala 12:21]
  assign _T_1537 = _T_1535 | _T_1536; // @[LZD.scala 49:16]
  assign _T_1538 = ~ _T_1536; // @[LZD.scala 49:27]
  assign _T_1539 = _T_1535 | _T_1538; // @[LZD.scala 49:25]
  assign _T_1540 = _T_1527[0:0]; // @[LZD.scala 49:47]
  assign _T_1541 = _T_1534[0:0]; // @[LZD.scala 49:59]
  assign _T_1542 = _T_1535 ? _T_1540 : _T_1541; // @[LZD.scala 49:35]
  assign _T_1544 = {_T_1537,_T_1539,_T_1542}; // @[Cat.scala 29:58]
  assign _T_1545 = _T_1519[2]; // @[Shift.scala 12:21]
  assign _T_1546 = _T_1544[2]; // @[Shift.scala 12:21]
  assign _T_1547 = _T_1545 | _T_1546; // @[LZD.scala 49:16]
  assign _T_1548 = ~ _T_1546; // @[LZD.scala 49:27]
  assign _T_1549 = _T_1545 | _T_1548; // @[LZD.scala 49:25]
  assign _T_1550 = _T_1519[1:0]; // @[LZD.scala 49:47]
  assign _T_1551 = _T_1544[1:0]; // @[LZD.scala 49:59]
  assign _T_1552 = _T_1545 ? _T_1550 : _T_1551; // @[LZD.scala 49:35]
  assign _T_1554 = {_T_1547,_T_1549,_T_1552}; // @[Cat.scala 29:58]
  assign _T_1555 = _T_1493[3]; // @[Shift.scala 12:21]
  assign _T_1556 = _T_1554[3]; // @[Shift.scala 12:21]
  assign _T_1557 = _T_1555 | _T_1556; // @[LZD.scala 49:16]
  assign _T_1558 = ~ _T_1556; // @[LZD.scala 49:27]
  assign _T_1559 = _T_1555 | _T_1558; // @[LZD.scala 49:25]
  assign _T_1560 = _T_1493[2:0]; // @[LZD.scala 49:47]
  assign _T_1561 = _T_1554[2:0]; // @[LZD.scala 49:59]
  assign _T_1562 = _T_1555 ? _T_1560 : _T_1561; // @[LZD.scala 49:35]
  assign _T_1564 = {_T_1557,_T_1559,_T_1562}; // @[Cat.scala 29:58]
  assign _T_1565 = _T_1431[15:0]; // @[LZD.scala 44:32]
  assign _T_1566 = _T_1565[15:8]; // @[LZD.scala 43:32]
  assign _T_1567 = _T_1566[7:4]; // @[LZD.scala 43:32]
  assign _T_1568 = _T_1567[3:2]; // @[LZD.scala 43:32]
  assign _T_1569 = _T_1568 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1570 = _T_1568[1]; // @[LZD.scala 39:21]
  assign _T_1571 = _T_1568[0]; // @[LZD.scala 39:30]
  assign _T_1572 = ~ _T_1571; // @[LZD.scala 39:27]
  assign _T_1573 = _T_1570 | _T_1572; // @[LZD.scala 39:25]
  assign _T_1574 = {_T_1569,_T_1573}; // @[Cat.scala 29:58]
  assign _T_1575 = _T_1567[1:0]; // @[LZD.scala 44:32]
  assign _T_1576 = _T_1575 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1577 = _T_1575[1]; // @[LZD.scala 39:21]
  assign _T_1578 = _T_1575[0]; // @[LZD.scala 39:30]
  assign _T_1579 = ~ _T_1578; // @[LZD.scala 39:27]
  assign _T_1580 = _T_1577 | _T_1579; // @[LZD.scala 39:25]
  assign _T_1581 = {_T_1576,_T_1580}; // @[Cat.scala 29:58]
  assign _T_1582 = _T_1574[1]; // @[Shift.scala 12:21]
  assign _T_1583 = _T_1581[1]; // @[Shift.scala 12:21]
  assign _T_1584 = _T_1582 | _T_1583; // @[LZD.scala 49:16]
  assign _T_1585 = ~ _T_1583; // @[LZD.scala 49:27]
  assign _T_1586 = _T_1582 | _T_1585; // @[LZD.scala 49:25]
  assign _T_1587 = _T_1574[0:0]; // @[LZD.scala 49:47]
  assign _T_1588 = _T_1581[0:0]; // @[LZD.scala 49:59]
  assign _T_1589 = _T_1582 ? _T_1587 : _T_1588; // @[LZD.scala 49:35]
  assign _T_1591 = {_T_1584,_T_1586,_T_1589}; // @[Cat.scala 29:58]
  assign _T_1592 = _T_1566[3:0]; // @[LZD.scala 44:32]
  assign _T_1593 = _T_1592[3:2]; // @[LZD.scala 43:32]
  assign _T_1594 = _T_1593 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1595 = _T_1593[1]; // @[LZD.scala 39:21]
  assign _T_1596 = _T_1593[0]; // @[LZD.scala 39:30]
  assign _T_1597 = ~ _T_1596; // @[LZD.scala 39:27]
  assign _T_1598 = _T_1595 | _T_1597; // @[LZD.scala 39:25]
  assign _T_1599 = {_T_1594,_T_1598}; // @[Cat.scala 29:58]
  assign _T_1600 = _T_1592[1:0]; // @[LZD.scala 44:32]
  assign _T_1601 = _T_1600 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1602 = _T_1600[1]; // @[LZD.scala 39:21]
  assign _T_1603 = _T_1600[0]; // @[LZD.scala 39:30]
  assign _T_1604 = ~ _T_1603; // @[LZD.scala 39:27]
  assign _T_1605 = _T_1602 | _T_1604; // @[LZD.scala 39:25]
  assign _T_1606 = {_T_1601,_T_1605}; // @[Cat.scala 29:58]
  assign _T_1607 = _T_1599[1]; // @[Shift.scala 12:21]
  assign _T_1608 = _T_1606[1]; // @[Shift.scala 12:21]
  assign _T_1609 = _T_1607 | _T_1608; // @[LZD.scala 49:16]
  assign _T_1610 = ~ _T_1608; // @[LZD.scala 49:27]
  assign _T_1611 = _T_1607 | _T_1610; // @[LZD.scala 49:25]
  assign _T_1612 = _T_1599[0:0]; // @[LZD.scala 49:47]
  assign _T_1613 = _T_1606[0:0]; // @[LZD.scala 49:59]
  assign _T_1614 = _T_1607 ? _T_1612 : _T_1613; // @[LZD.scala 49:35]
  assign _T_1616 = {_T_1609,_T_1611,_T_1614}; // @[Cat.scala 29:58]
  assign _T_1617 = _T_1591[2]; // @[Shift.scala 12:21]
  assign _T_1618 = _T_1616[2]; // @[Shift.scala 12:21]
  assign _T_1619 = _T_1617 | _T_1618; // @[LZD.scala 49:16]
  assign _T_1620 = ~ _T_1618; // @[LZD.scala 49:27]
  assign _T_1621 = _T_1617 | _T_1620; // @[LZD.scala 49:25]
  assign _T_1622 = _T_1591[1:0]; // @[LZD.scala 49:47]
  assign _T_1623 = _T_1616[1:0]; // @[LZD.scala 49:59]
  assign _T_1624 = _T_1617 ? _T_1622 : _T_1623; // @[LZD.scala 49:35]
  assign _T_1626 = {_T_1619,_T_1621,_T_1624}; // @[Cat.scala 29:58]
  assign _T_1627 = _T_1565[7:0]; // @[LZD.scala 44:32]
  assign _T_1628 = _T_1627[7:4]; // @[LZD.scala 43:32]
  assign _T_1629 = _T_1628[3:2]; // @[LZD.scala 43:32]
  assign _T_1630 = _T_1629 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1631 = _T_1629[1]; // @[LZD.scala 39:21]
  assign _T_1632 = _T_1629[0]; // @[LZD.scala 39:30]
  assign _T_1633 = ~ _T_1632; // @[LZD.scala 39:27]
  assign _T_1634 = _T_1631 | _T_1633; // @[LZD.scala 39:25]
  assign _T_1635 = {_T_1630,_T_1634}; // @[Cat.scala 29:58]
  assign _T_1636 = _T_1628[1:0]; // @[LZD.scala 44:32]
  assign _T_1637 = _T_1636 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1638 = _T_1636[1]; // @[LZD.scala 39:21]
  assign _T_1639 = _T_1636[0]; // @[LZD.scala 39:30]
  assign _T_1640 = ~ _T_1639; // @[LZD.scala 39:27]
  assign _T_1641 = _T_1638 | _T_1640; // @[LZD.scala 39:25]
  assign _T_1642 = {_T_1637,_T_1641}; // @[Cat.scala 29:58]
  assign _T_1643 = _T_1635[1]; // @[Shift.scala 12:21]
  assign _T_1644 = _T_1642[1]; // @[Shift.scala 12:21]
  assign _T_1645 = _T_1643 | _T_1644; // @[LZD.scala 49:16]
  assign _T_1646 = ~ _T_1644; // @[LZD.scala 49:27]
  assign _T_1647 = _T_1643 | _T_1646; // @[LZD.scala 49:25]
  assign _T_1648 = _T_1635[0:0]; // @[LZD.scala 49:47]
  assign _T_1649 = _T_1642[0:0]; // @[LZD.scala 49:59]
  assign _T_1650 = _T_1643 ? _T_1648 : _T_1649; // @[LZD.scala 49:35]
  assign _T_1652 = {_T_1645,_T_1647,_T_1650}; // @[Cat.scala 29:58]
  assign _T_1653 = _T_1627[3:0]; // @[LZD.scala 44:32]
  assign _T_1654 = _T_1653[3:2]; // @[LZD.scala 43:32]
  assign _T_1655 = _T_1654 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1656 = _T_1654[1]; // @[LZD.scala 39:21]
  assign _T_1657 = _T_1654[0]; // @[LZD.scala 39:30]
  assign _T_1658 = ~ _T_1657; // @[LZD.scala 39:27]
  assign _T_1659 = _T_1656 | _T_1658; // @[LZD.scala 39:25]
  assign _T_1660 = {_T_1655,_T_1659}; // @[Cat.scala 29:58]
  assign _T_1661 = _T_1653[1:0]; // @[LZD.scala 44:32]
  assign _T_1662 = _T_1661 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1663 = _T_1661[1]; // @[LZD.scala 39:21]
  assign _T_1664 = _T_1661[0]; // @[LZD.scala 39:30]
  assign _T_1665 = ~ _T_1664; // @[LZD.scala 39:27]
  assign _T_1666 = _T_1663 | _T_1665; // @[LZD.scala 39:25]
  assign _T_1667 = {_T_1662,_T_1666}; // @[Cat.scala 29:58]
  assign _T_1668 = _T_1660[1]; // @[Shift.scala 12:21]
  assign _T_1669 = _T_1667[1]; // @[Shift.scala 12:21]
  assign _T_1670 = _T_1668 | _T_1669; // @[LZD.scala 49:16]
  assign _T_1671 = ~ _T_1669; // @[LZD.scala 49:27]
  assign _T_1672 = _T_1668 | _T_1671; // @[LZD.scala 49:25]
  assign _T_1673 = _T_1660[0:0]; // @[LZD.scala 49:47]
  assign _T_1674 = _T_1667[0:0]; // @[LZD.scala 49:59]
  assign _T_1675 = _T_1668 ? _T_1673 : _T_1674; // @[LZD.scala 49:35]
  assign _T_1677 = {_T_1670,_T_1672,_T_1675}; // @[Cat.scala 29:58]
  assign _T_1678 = _T_1652[2]; // @[Shift.scala 12:21]
  assign _T_1679 = _T_1677[2]; // @[Shift.scala 12:21]
  assign _T_1680 = _T_1678 | _T_1679; // @[LZD.scala 49:16]
  assign _T_1681 = ~ _T_1679; // @[LZD.scala 49:27]
  assign _T_1682 = _T_1678 | _T_1681; // @[LZD.scala 49:25]
  assign _T_1683 = _T_1652[1:0]; // @[LZD.scala 49:47]
  assign _T_1684 = _T_1677[1:0]; // @[LZD.scala 49:59]
  assign _T_1685 = _T_1678 ? _T_1683 : _T_1684; // @[LZD.scala 49:35]
  assign _T_1687 = {_T_1680,_T_1682,_T_1685}; // @[Cat.scala 29:58]
  assign _T_1688 = _T_1626[3]; // @[Shift.scala 12:21]
  assign _T_1689 = _T_1687[3]; // @[Shift.scala 12:21]
  assign _T_1690 = _T_1688 | _T_1689; // @[LZD.scala 49:16]
  assign _T_1691 = ~ _T_1689; // @[LZD.scala 49:27]
  assign _T_1692 = _T_1688 | _T_1691; // @[LZD.scala 49:25]
  assign _T_1693 = _T_1626[2:0]; // @[LZD.scala 49:47]
  assign _T_1694 = _T_1687[2:0]; // @[LZD.scala 49:59]
  assign _T_1695 = _T_1688 ? _T_1693 : _T_1694; // @[LZD.scala 49:35]
  assign _T_1697 = {_T_1690,_T_1692,_T_1695}; // @[Cat.scala 29:58]
  assign _T_1698 = _T_1564[4]; // @[Shift.scala 12:21]
  assign _T_1699 = _T_1697[4]; // @[Shift.scala 12:21]
  assign _T_1700 = _T_1698 | _T_1699; // @[LZD.scala 49:16]
  assign _T_1701 = ~ _T_1699; // @[LZD.scala 49:27]
  assign _T_1702 = _T_1698 | _T_1701; // @[LZD.scala 49:25]
  assign _T_1703 = _T_1564[3:0]; // @[LZD.scala 49:47]
  assign _T_1704 = _T_1697[3:0]; // @[LZD.scala 49:59]
  assign _T_1705 = _T_1698 ? _T_1703 : _T_1704; // @[LZD.scala 49:35]
  assign _T_1707 = {_T_1700,_T_1702,_T_1705}; // @[Cat.scala 29:58]
  assign _T_1708 = _T_1430[5]; // @[Shift.scala 12:21]
  assign _T_1709 = _T_1707[5]; // @[Shift.scala 12:21]
  assign _T_1710 = _T_1708 | _T_1709; // @[LZD.scala 49:16]
  assign _T_1711 = ~ _T_1709; // @[LZD.scala 49:27]
  assign _T_1712 = _T_1708 | _T_1711; // @[LZD.scala 49:25]
  assign _T_1713 = _T_1430[4:0]; // @[LZD.scala 49:47]
  assign _T_1714 = _T_1707[4:0]; // @[LZD.scala 49:59]
  assign _T_1715 = _T_1708 ? _T_1713 : _T_1714; // @[LZD.scala 49:35]
  assign _T_1717 = {_T_1710,_T_1712,_T_1715}; // @[Cat.scala 29:58]
  assign _T_1718 = _T_1152[63:0]; // @[LZD.scala 44:32]
  assign _T_1719 = _T_1718[63:32]; // @[LZD.scala 43:32]
  assign _T_1720 = _T_1719[31:16]; // @[LZD.scala 43:32]
  assign _T_1721 = _T_1720[15:8]; // @[LZD.scala 43:32]
  assign _T_1722 = _T_1721[7:4]; // @[LZD.scala 43:32]
  assign _T_1723 = _T_1722[3:2]; // @[LZD.scala 43:32]
  assign _T_1724 = _T_1723 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1725 = _T_1723[1]; // @[LZD.scala 39:21]
  assign _T_1726 = _T_1723[0]; // @[LZD.scala 39:30]
  assign _T_1727 = ~ _T_1726; // @[LZD.scala 39:27]
  assign _T_1728 = _T_1725 | _T_1727; // @[LZD.scala 39:25]
  assign _T_1729 = {_T_1724,_T_1728}; // @[Cat.scala 29:58]
  assign _T_1730 = _T_1722[1:0]; // @[LZD.scala 44:32]
  assign _T_1731 = _T_1730 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1732 = _T_1730[1]; // @[LZD.scala 39:21]
  assign _T_1733 = _T_1730[0]; // @[LZD.scala 39:30]
  assign _T_1734 = ~ _T_1733; // @[LZD.scala 39:27]
  assign _T_1735 = _T_1732 | _T_1734; // @[LZD.scala 39:25]
  assign _T_1736 = {_T_1731,_T_1735}; // @[Cat.scala 29:58]
  assign _T_1737 = _T_1729[1]; // @[Shift.scala 12:21]
  assign _T_1738 = _T_1736[1]; // @[Shift.scala 12:21]
  assign _T_1739 = _T_1737 | _T_1738; // @[LZD.scala 49:16]
  assign _T_1740 = ~ _T_1738; // @[LZD.scala 49:27]
  assign _T_1741 = _T_1737 | _T_1740; // @[LZD.scala 49:25]
  assign _T_1742 = _T_1729[0:0]; // @[LZD.scala 49:47]
  assign _T_1743 = _T_1736[0:0]; // @[LZD.scala 49:59]
  assign _T_1744 = _T_1737 ? _T_1742 : _T_1743; // @[LZD.scala 49:35]
  assign _T_1746 = {_T_1739,_T_1741,_T_1744}; // @[Cat.scala 29:58]
  assign _T_1747 = _T_1721[3:0]; // @[LZD.scala 44:32]
  assign _T_1748 = _T_1747[3:2]; // @[LZD.scala 43:32]
  assign _T_1749 = _T_1748 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1750 = _T_1748[1]; // @[LZD.scala 39:21]
  assign _T_1751 = _T_1748[0]; // @[LZD.scala 39:30]
  assign _T_1752 = ~ _T_1751; // @[LZD.scala 39:27]
  assign _T_1753 = _T_1750 | _T_1752; // @[LZD.scala 39:25]
  assign _T_1754 = {_T_1749,_T_1753}; // @[Cat.scala 29:58]
  assign _T_1755 = _T_1747[1:0]; // @[LZD.scala 44:32]
  assign _T_1756 = _T_1755 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1757 = _T_1755[1]; // @[LZD.scala 39:21]
  assign _T_1758 = _T_1755[0]; // @[LZD.scala 39:30]
  assign _T_1759 = ~ _T_1758; // @[LZD.scala 39:27]
  assign _T_1760 = _T_1757 | _T_1759; // @[LZD.scala 39:25]
  assign _T_1761 = {_T_1756,_T_1760}; // @[Cat.scala 29:58]
  assign _T_1762 = _T_1754[1]; // @[Shift.scala 12:21]
  assign _T_1763 = _T_1761[1]; // @[Shift.scala 12:21]
  assign _T_1764 = _T_1762 | _T_1763; // @[LZD.scala 49:16]
  assign _T_1765 = ~ _T_1763; // @[LZD.scala 49:27]
  assign _T_1766 = _T_1762 | _T_1765; // @[LZD.scala 49:25]
  assign _T_1767 = _T_1754[0:0]; // @[LZD.scala 49:47]
  assign _T_1768 = _T_1761[0:0]; // @[LZD.scala 49:59]
  assign _T_1769 = _T_1762 ? _T_1767 : _T_1768; // @[LZD.scala 49:35]
  assign _T_1771 = {_T_1764,_T_1766,_T_1769}; // @[Cat.scala 29:58]
  assign _T_1772 = _T_1746[2]; // @[Shift.scala 12:21]
  assign _T_1773 = _T_1771[2]; // @[Shift.scala 12:21]
  assign _T_1774 = _T_1772 | _T_1773; // @[LZD.scala 49:16]
  assign _T_1775 = ~ _T_1773; // @[LZD.scala 49:27]
  assign _T_1776 = _T_1772 | _T_1775; // @[LZD.scala 49:25]
  assign _T_1777 = _T_1746[1:0]; // @[LZD.scala 49:47]
  assign _T_1778 = _T_1771[1:0]; // @[LZD.scala 49:59]
  assign _T_1779 = _T_1772 ? _T_1777 : _T_1778; // @[LZD.scala 49:35]
  assign _T_1781 = {_T_1774,_T_1776,_T_1779}; // @[Cat.scala 29:58]
  assign _T_1782 = _T_1720[7:0]; // @[LZD.scala 44:32]
  assign _T_1783 = _T_1782[7:4]; // @[LZD.scala 43:32]
  assign _T_1784 = _T_1783[3:2]; // @[LZD.scala 43:32]
  assign _T_1785 = _T_1784 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1786 = _T_1784[1]; // @[LZD.scala 39:21]
  assign _T_1787 = _T_1784[0]; // @[LZD.scala 39:30]
  assign _T_1788 = ~ _T_1787; // @[LZD.scala 39:27]
  assign _T_1789 = _T_1786 | _T_1788; // @[LZD.scala 39:25]
  assign _T_1790 = {_T_1785,_T_1789}; // @[Cat.scala 29:58]
  assign _T_1791 = _T_1783[1:0]; // @[LZD.scala 44:32]
  assign _T_1792 = _T_1791 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1793 = _T_1791[1]; // @[LZD.scala 39:21]
  assign _T_1794 = _T_1791[0]; // @[LZD.scala 39:30]
  assign _T_1795 = ~ _T_1794; // @[LZD.scala 39:27]
  assign _T_1796 = _T_1793 | _T_1795; // @[LZD.scala 39:25]
  assign _T_1797 = {_T_1792,_T_1796}; // @[Cat.scala 29:58]
  assign _T_1798 = _T_1790[1]; // @[Shift.scala 12:21]
  assign _T_1799 = _T_1797[1]; // @[Shift.scala 12:21]
  assign _T_1800 = _T_1798 | _T_1799; // @[LZD.scala 49:16]
  assign _T_1801 = ~ _T_1799; // @[LZD.scala 49:27]
  assign _T_1802 = _T_1798 | _T_1801; // @[LZD.scala 49:25]
  assign _T_1803 = _T_1790[0:0]; // @[LZD.scala 49:47]
  assign _T_1804 = _T_1797[0:0]; // @[LZD.scala 49:59]
  assign _T_1805 = _T_1798 ? _T_1803 : _T_1804; // @[LZD.scala 49:35]
  assign _T_1807 = {_T_1800,_T_1802,_T_1805}; // @[Cat.scala 29:58]
  assign _T_1808 = _T_1782[3:0]; // @[LZD.scala 44:32]
  assign _T_1809 = _T_1808[3:2]; // @[LZD.scala 43:32]
  assign _T_1810 = _T_1809 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1811 = _T_1809[1]; // @[LZD.scala 39:21]
  assign _T_1812 = _T_1809[0]; // @[LZD.scala 39:30]
  assign _T_1813 = ~ _T_1812; // @[LZD.scala 39:27]
  assign _T_1814 = _T_1811 | _T_1813; // @[LZD.scala 39:25]
  assign _T_1815 = {_T_1810,_T_1814}; // @[Cat.scala 29:58]
  assign _T_1816 = _T_1808[1:0]; // @[LZD.scala 44:32]
  assign _T_1817 = _T_1816 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1818 = _T_1816[1]; // @[LZD.scala 39:21]
  assign _T_1819 = _T_1816[0]; // @[LZD.scala 39:30]
  assign _T_1820 = ~ _T_1819; // @[LZD.scala 39:27]
  assign _T_1821 = _T_1818 | _T_1820; // @[LZD.scala 39:25]
  assign _T_1822 = {_T_1817,_T_1821}; // @[Cat.scala 29:58]
  assign _T_1823 = _T_1815[1]; // @[Shift.scala 12:21]
  assign _T_1824 = _T_1822[1]; // @[Shift.scala 12:21]
  assign _T_1825 = _T_1823 | _T_1824; // @[LZD.scala 49:16]
  assign _T_1826 = ~ _T_1824; // @[LZD.scala 49:27]
  assign _T_1827 = _T_1823 | _T_1826; // @[LZD.scala 49:25]
  assign _T_1828 = _T_1815[0:0]; // @[LZD.scala 49:47]
  assign _T_1829 = _T_1822[0:0]; // @[LZD.scala 49:59]
  assign _T_1830 = _T_1823 ? _T_1828 : _T_1829; // @[LZD.scala 49:35]
  assign _T_1832 = {_T_1825,_T_1827,_T_1830}; // @[Cat.scala 29:58]
  assign _T_1833 = _T_1807[2]; // @[Shift.scala 12:21]
  assign _T_1834 = _T_1832[2]; // @[Shift.scala 12:21]
  assign _T_1835 = _T_1833 | _T_1834; // @[LZD.scala 49:16]
  assign _T_1836 = ~ _T_1834; // @[LZD.scala 49:27]
  assign _T_1837 = _T_1833 | _T_1836; // @[LZD.scala 49:25]
  assign _T_1838 = _T_1807[1:0]; // @[LZD.scala 49:47]
  assign _T_1839 = _T_1832[1:0]; // @[LZD.scala 49:59]
  assign _T_1840 = _T_1833 ? _T_1838 : _T_1839; // @[LZD.scala 49:35]
  assign _T_1842 = {_T_1835,_T_1837,_T_1840}; // @[Cat.scala 29:58]
  assign _T_1843 = _T_1781[3]; // @[Shift.scala 12:21]
  assign _T_1844 = _T_1842[3]; // @[Shift.scala 12:21]
  assign _T_1845 = _T_1843 | _T_1844; // @[LZD.scala 49:16]
  assign _T_1846 = ~ _T_1844; // @[LZD.scala 49:27]
  assign _T_1847 = _T_1843 | _T_1846; // @[LZD.scala 49:25]
  assign _T_1848 = _T_1781[2:0]; // @[LZD.scala 49:47]
  assign _T_1849 = _T_1842[2:0]; // @[LZD.scala 49:59]
  assign _T_1850 = _T_1843 ? _T_1848 : _T_1849; // @[LZD.scala 49:35]
  assign _T_1852 = {_T_1845,_T_1847,_T_1850}; // @[Cat.scala 29:58]
  assign _T_1853 = _T_1719[15:0]; // @[LZD.scala 44:32]
  assign _T_1854 = _T_1853[15:8]; // @[LZD.scala 43:32]
  assign _T_1855 = _T_1854[7:4]; // @[LZD.scala 43:32]
  assign _T_1856 = _T_1855[3:2]; // @[LZD.scala 43:32]
  assign _T_1857 = _T_1856 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1858 = _T_1856[1]; // @[LZD.scala 39:21]
  assign _T_1859 = _T_1856[0]; // @[LZD.scala 39:30]
  assign _T_1860 = ~ _T_1859; // @[LZD.scala 39:27]
  assign _T_1861 = _T_1858 | _T_1860; // @[LZD.scala 39:25]
  assign _T_1862 = {_T_1857,_T_1861}; // @[Cat.scala 29:58]
  assign _T_1863 = _T_1855[1:0]; // @[LZD.scala 44:32]
  assign _T_1864 = _T_1863 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1865 = _T_1863[1]; // @[LZD.scala 39:21]
  assign _T_1866 = _T_1863[0]; // @[LZD.scala 39:30]
  assign _T_1867 = ~ _T_1866; // @[LZD.scala 39:27]
  assign _T_1868 = _T_1865 | _T_1867; // @[LZD.scala 39:25]
  assign _T_1869 = {_T_1864,_T_1868}; // @[Cat.scala 29:58]
  assign _T_1870 = _T_1862[1]; // @[Shift.scala 12:21]
  assign _T_1871 = _T_1869[1]; // @[Shift.scala 12:21]
  assign _T_1872 = _T_1870 | _T_1871; // @[LZD.scala 49:16]
  assign _T_1873 = ~ _T_1871; // @[LZD.scala 49:27]
  assign _T_1874 = _T_1870 | _T_1873; // @[LZD.scala 49:25]
  assign _T_1875 = _T_1862[0:0]; // @[LZD.scala 49:47]
  assign _T_1876 = _T_1869[0:0]; // @[LZD.scala 49:59]
  assign _T_1877 = _T_1870 ? _T_1875 : _T_1876; // @[LZD.scala 49:35]
  assign _T_1879 = {_T_1872,_T_1874,_T_1877}; // @[Cat.scala 29:58]
  assign _T_1880 = _T_1854[3:0]; // @[LZD.scala 44:32]
  assign _T_1881 = _T_1880[3:2]; // @[LZD.scala 43:32]
  assign _T_1882 = _T_1881 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1883 = _T_1881[1]; // @[LZD.scala 39:21]
  assign _T_1884 = _T_1881[0]; // @[LZD.scala 39:30]
  assign _T_1885 = ~ _T_1884; // @[LZD.scala 39:27]
  assign _T_1886 = _T_1883 | _T_1885; // @[LZD.scala 39:25]
  assign _T_1887 = {_T_1882,_T_1886}; // @[Cat.scala 29:58]
  assign _T_1888 = _T_1880[1:0]; // @[LZD.scala 44:32]
  assign _T_1889 = _T_1888 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1890 = _T_1888[1]; // @[LZD.scala 39:21]
  assign _T_1891 = _T_1888[0]; // @[LZD.scala 39:30]
  assign _T_1892 = ~ _T_1891; // @[LZD.scala 39:27]
  assign _T_1893 = _T_1890 | _T_1892; // @[LZD.scala 39:25]
  assign _T_1894 = {_T_1889,_T_1893}; // @[Cat.scala 29:58]
  assign _T_1895 = _T_1887[1]; // @[Shift.scala 12:21]
  assign _T_1896 = _T_1894[1]; // @[Shift.scala 12:21]
  assign _T_1897 = _T_1895 | _T_1896; // @[LZD.scala 49:16]
  assign _T_1898 = ~ _T_1896; // @[LZD.scala 49:27]
  assign _T_1899 = _T_1895 | _T_1898; // @[LZD.scala 49:25]
  assign _T_1900 = _T_1887[0:0]; // @[LZD.scala 49:47]
  assign _T_1901 = _T_1894[0:0]; // @[LZD.scala 49:59]
  assign _T_1902 = _T_1895 ? _T_1900 : _T_1901; // @[LZD.scala 49:35]
  assign _T_1904 = {_T_1897,_T_1899,_T_1902}; // @[Cat.scala 29:58]
  assign _T_1905 = _T_1879[2]; // @[Shift.scala 12:21]
  assign _T_1906 = _T_1904[2]; // @[Shift.scala 12:21]
  assign _T_1907 = _T_1905 | _T_1906; // @[LZD.scala 49:16]
  assign _T_1908 = ~ _T_1906; // @[LZD.scala 49:27]
  assign _T_1909 = _T_1905 | _T_1908; // @[LZD.scala 49:25]
  assign _T_1910 = _T_1879[1:0]; // @[LZD.scala 49:47]
  assign _T_1911 = _T_1904[1:0]; // @[LZD.scala 49:59]
  assign _T_1912 = _T_1905 ? _T_1910 : _T_1911; // @[LZD.scala 49:35]
  assign _T_1914 = {_T_1907,_T_1909,_T_1912}; // @[Cat.scala 29:58]
  assign _T_1915 = _T_1853[7:0]; // @[LZD.scala 44:32]
  assign _T_1916 = _T_1915[7:4]; // @[LZD.scala 43:32]
  assign _T_1917 = _T_1916[3:2]; // @[LZD.scala 43:32]
  assign _T_1918 = _T_1917 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1919 = _T_1917[1]; // @[LZD.scala 39:21]
  assign _T_1920 = _T_1917[0]; // @[LZD.scala 39:30]
  assign _T_1921 = ~ _T_1920; // @[LZD.scala 39:27]
  assign _T_1922 = _T_1919 | _T_1921; // @[LZD.scala 39:25]
  assign _T_1923 = {_T_1918,_T_1922}; // @[Cat.scala 29:58]
  assign _T_1924 = _T_1916[1:0]; // @[LZD.scala 44:32]
  assign _T_1925 = _T_1924 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1926 = _T_1924[1]; // @[LZD.scala 39:21]
  assign _T_1927 = _T_1924[0]; // @[LZD.scala 39:30]
  assign _T_1928 = ~ _T_1927; // @[LZD.scala 39:27]
  assign _T_1929 = _T_1926 | _T_1928; // @[LZD.scala 39:25]
  assign _T_1930 = {_T_1925,_T_1929}; // @[Cat.scala 29:58]
  assign _T_1931 = _T_1923[1]; // @[Shift.scala 12:21]
  assign _T_1932 = _T_1930[1]; // @[Shift.scala 12:21]
  assign _T_1933 = _T_1931 | _T_1932; // @[LZD.scala 49:16]
  assign _T_1934 = ~ _T_1932; // @[LZD.scala 49:27]
  assign _T_1935 = _T_1931 | _T_1934; // @[LZD.scala 49:25]
  assign _T_1936 = _T_1923[0:0]; // @[LZD.scala 49:47]
  assign _T_1937 = _T_1930[0:0]; // @[LZD.scala 49:59]
  assign _T_1938 = _T_1931 ? _T_1936 : _T_1937; // @[LZD.scala 49:35]
  assign _T_1940 = {_T_1933,_T_1935,_T_1938}; // @[Cat.scala 29:58]
  assign _T_1941 = _T_1915[3:0]; // @[LZD.scala 44:32]
  assign _T_1942 = _T_1941[3:2]; // @[LZD.scala 43:32]
  assign _T_1943 = _T_1942 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1944 = _T_1942[1]; // @[LZD.scala 39:21]
  assign _T_1945 = _T_1942[0]; // @[LZD.scala 39:30]
  assign _T_1946 = ~ _T_1945; // @[LZD.scala 39:27]
  assign _T_1947 = _T_1944 | _T_1946; // @[LZD.scala 39:25]
  assign _T_1948 = {_T_1943,_T_1947}; // @[Cat.scala 29:58]
  assign _T_1949 = _T_1941[1:0]; // @[LZD.scala 44:32]
  assign _T_1950 = _T_1949 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1951 = _T_1949[1]; // @[LZD.scala 39:21]
  assign _T_1952 = _T_1949[0]; // @[LZD.scala 39:30]
  assign _T_1953 = ~ _T_1952; // @[LZD.scala 39:27]
  assign _T_1954 = _T_1951 | _T_1953; // @[LZD.scala 39:25]
  assign _T_1955 = {_T_1950,_T_1954}; // @[Cat.scala 29:58]
  assign _T_1956 = _T_1948[1]; // @[Shift.scala 12:21]
  assign _T_1957 = _T_1955[1]; // @[Shift.scala 12:21]
  assign _T_1958 = _T_1956 | _T_1957; // @[LZD.scala 49:16]
  assign _T_1959 = ~ _T_1957; // @[LZD.scala 49:27]
  assign _T_1960 = _T_1956 | _T_1959; // @[LZD.scala 49:25]
  assign _T_1961 = _T_1948[0:0]; // @[LZD.scala 49:47]
  assign _T_1962 = _T_1955[0:0]; // @[LZD.scala 49:59]
  assign _T_1963 = _T_1956 ? _T_1961 : _T_1962; // @[LZD.scala 49:35]
  assign _T_1965 = {_T_1958,_T_1960,_T_1963}; // @[Cat.scala 29:58]
  assign _T_1966 = _T_1940[2]; // @[Shift.scala 12:21]
  assign _T_1967 = _T_1965[2]; // @[Shift.scala 12:21]
  assign _T_1968 = _T_1966 | _T_1967; // @[LZD.scala 49:16]
  assign _T_1969 = ~ _T_1967; // @[LZD.scala 49:27]
  assign _T_1970 = _T_1966 | _T_1969; // @[LZD.scala 49:25]
  assign _T_1971 = _T_1940[1:0]; // @[LZD.scala 49:47]
  assign _T_1972 = _T_1965[1:0]; // @[LZD.scala 49:59]
  assign _T_1973 = _T_1966 ? _T_1971 : _T_1972; // @[LZD.scala 49:35]
  assign _T_1975 = {_T_1968,_T_1970,_T_1973}; // @[Cat.scala 29:58]
  assign _T_1976 = _T_1914[3]; // @[Shift.scala 12:21]
  assign _T_1977 = _T_1975[3]; // @[Shift.scala 12:21]
  assign _T_1978 = _T_1976 | _T_1977; // @[LZD.scala 49:16]
  assign _T_1979 = ~ _T_1977; // @[LZD.scala 49:27]
  assign _T_1980 = _T_1976 | _T_1979; // @[LZD.scala 49:25]
  assign _T_1981 = _T_1914[2:0]; // @[LZD.scala 49:47]
  assign _T_1982 = _T_1975[2:0]; // @[LZD.scala 49:59]
  assign _T_1983 = _T_1976 ? _T_1981 : _T_1982; // @[LZD.scala 49:35]
  assign _T_1985 = {_T_1978,_T_1980,_T_1983}; // @[Cat.scala 29:58]
  assign _T_1986 = _T_1852[4]; // @[Shift.scala 12:21]
  assign _T_1987 = _T_1985[4]; // @[Shift.scala 12:21]
  assign _T_1988 = _T_1986 | _T_1987; // @[LZD.scala 49:16]
  assign _T_1989 = ~ _T_1987; // @[LZD.scala 49:27]
  assign _T_1990 = _T_1986 | _T_1989; // @[LZD.scala 49:25]
  assign _T_1991 = _T_1852[3:0]; // @[LZD.scala 49:47]
  assign _T_1992 = _T_1985[3:0]; // @[LZD.scala 49:59]
  assign _T_1993 = _T_1986 ? _T_1991 : _T_1992; // @[LZD.scala 49:35]
  assign _T_1995 = {_T_1988,_T_1990,_T_1993}; // @[Cat.scala 29:58]
  assign _T_1996 = _T_1718[31:0]; // @[LZD.scala 44:32]
  assign _T_1997 = _T_1996[31:16]; // @[LZD.scala 43:32]
  assign _T_1998 = _T_1997[15:8]; // @[LZD.scala 43:32]
  assign _T_1999 = _T_1998[7:4]; // @[LZD.scala 43:32]
  assign _T_2000 = _T_1999[3:2]; // @[LZD.scala 43:32]
  assign _T_2001 = _T_2000 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2002 = _T_2000[1]; // @[LZD.scala 39:21]
  assign _T_2003 = _T_2000[0]; // @[LZD.scala 39:30]
  assign _T_2004 = ~ _T_2003; // @[LZD.scala 39:27]
  assign _T_2005 = _T_2002 | _T_2004; // @[LZD.scala 39:25]
  assign _T_2006 = {_T_2001,_T_2005}; // @[Cat.scala 29:58]
  assign _T_2007 = _T_1999[1:0]; // @[LZD.scala 44:32]
  assign _T_2008 = _T_2007 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2009 = _T_2007[1]; // @[LZD.scala 39:21]
  assign _T_2010 = _T_2007[0]; // @[LZD.scala 39:30]
  assign _T_2011 = ~ _T_2010; // @[LZD.scala 39:27]
  assign _T_2012 = _T_2009 | _T_2011; // @[LZD.scala 39:25]
  assign _T_2013 = {_T_2008,_T_2012}; // @[Cat.scala 29:58]
  assign _T_2014 = _T_2006[1]; // @[Shift.scala 12:21]
  assign _T_2015 = _T_2013[1]; // @[Shift.scala 12:21]
  assign _T_2016 = _T_2014 | _T_2015; // @[LZD.scala 49:16]
  assign _T_2017 = ~ _T_2015; // @[LZD.scala 49:27]
  assign _T_2018 = _T_2014 | _T_2017; // @[LZD.scala 49:25]
  assign _T_2019 = _T_2006[0:0]; // @[LZD.scala 49:47]
  assign _T_2020 = _T_2013[0:0]; // @[LZD.scala 49:59]
  assign _T_2021 = _T_2014 ? _T_2019 : _T_2020; // @[LZD.scala 49:35]
  assign _T_2023 = {_T_2016,_T_2018,_T_2021}; // @[Cat.scala 29:58]
  assign _T_2024 = _T_1998[3:0]; // @[LZD.scala 44:32]
  assign _T_2025 = _T_2024[3:2]; // @[LZD.scala 43:32]
  assign _T_2026 = _T_2025 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2027 = _T_2025[1]; // @[LZD.scala 39:21]
  assign _T_2028 = _T_2025[0]; // @[LZD.scala 39:30]
  assign _T_2029 = ~ _T_2028; // @[LZD.scala 39:27]
  assign _T_2030 = _T_2027 | _T_2029; // @[LZD.scala 39:25]
  assign _T_2031 = {_T_2026,_T_2030}; // @[Cat.scala 29:58]
  assign _T_2032 = _T_2024[1:0]; // @[LZD.scala 44:32]
  assign _T_2033 = _T_2032 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2034 = _T_2032[1]; // @[LZD.scala 39:21]
  assign _T_2035 = _T_2032[0]; // @[LZD.scala 39:30]
  assign _T_2036 = ~ _T_2035; // @[LZD.scala 39:27]
  assign _T_2037 = _T_2034 | _T_2036; // @[LZD.scala 39:25]
  assign _T_2038 = {_T_2033,_T_2037}; // @[Cat.scala 29:58]
  assign _T_2039 = _T_2031[1]; // @[Shift.scala 12:21]
  assign _T_2040 = _T_2038[1]; // @[Shift.scala 12:21]
  assign _T_2041 = _T_2039 | _T_2040; // @[LZD.scala 49:16]
  assign _T_2042 = ~ _T_2040; // @[LZD.scala 49:27]
  assign _T_2043 = _T_2039 | _T_2042; // @[LZD.scala 49:25]
  assign _T_2044 = _T_2031[0:0]; // @[LZD.scala 49:47]
  assign _T_2045 = _T_2038[0:0]; // @[LZD.scala 49:59]
  assign _T_2046 = _T_2039 ? _T_2044 : _T_2045; // @[LZD.scala 49:35]
  assign _T_2048 = {_T_2041,_T_2043,_T_2046}; // @[Cat.scala 29:58]
  assign _T_2049 = _T_2023[2]; // @[Shift.scala 12:21]
  assign _T_2050 = _T_2048[2]; // @[Shift.scala 12:21]
  assign _T_2051 = _T_2049 | _T_2050; // @[LZD.scala 49:16]
  assign _T_2052 = ~ _T_2050; // @[LZD.scala 49:27]
  assign _T_2053 = _T_2049 | _T_2052; // @[LZD.scala 49:25]
  assign _T_2054 = _T_2023[1:0]; // @[LZD.scala 49:47]
  assign _T_2055 = _T_2048[1:0]; // @[LZD.scala 49:59]
  assign _T_2056 = _T_2049 ? _T_2054 : _T_2055; // @[LZD.scala 49:35]
  assign _T_2058 = {_T_2051,_T_2053,_T_2056}; // @[Cat.scala 29:58]
  assign _T_2059 = _T_1997[7:0]; // @[LZD.scala 44:32]
  assign _T_2060 = _T_2059[7:4]; // @[LZD.scala 43:32]
  assign _T_2061 = _T_2060[3:2]; // @[LZD.scala 43:32]
  assign _T_2062 = _T_2061 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2063 = _T_2061[1]; // @[LZD.scala 39:21]
  assign _T_2064 = _T_2061[0]; // @[LZD.scala 39:30]
  assign _T_2065 = ~ _T_2064; // @[LZD.scala 39:27]
  assign _T_2066 = _T_2063 | _T_2065; // @[LZD.scala 39:25]
  assign _T_2067 = {_T_2062,_T_2066}; // @[Cat.scala 29:58]
  assign _T_2068 = _T_2060[1:0]; // @[LZD.scala 44:32]
  assign _T_2069 = _T_2068 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2070 = _T_2068[1]; // @[LZD.scala 39:21]
  assign _T_2071 = _T_2068[0]; // @[LZD.scala 39:30]
  assign _T_2072 = ~ _T_2071; // @[LZD.scala 39:27]
  assign _T_2073 = _T_2070 | _T_2072; // @[LZD.scala 39:25]
  assign _T_2074 = {_T_2069,_T_2073}; // @[Cat.scala 29:58]
  assign _T_2075 = _T_2067[1]; // @[Shift.scala 12:21]
  assign _T_2076 = _T_2074[1]; // @[Shift.scala 12:21]
  assign _T_2077 = _T_2075 | _T_2076; // @[LZD.scala 49:16]
  assign _T_2078 = ~ _T_2076; // @[LZD.scala 49:27]
  assign _T_2079 = _T_2075 | _T_2078; // @[LZD.scala 49:25]
  assign _T_2080 = _T_2067[0:0]; // @[LZD.scala 49:47]
  assign _T_2081 = _T_2074[0:0]; // @[LZD.scala 49:59]
  assign _T_2082 = _T_2075 ? _T_2080 : _T_2081; // @[LZD.scala 49:35]
  assign _T_2084 = {_T_2077,_T_2079,_T_2082}; // @[Cat.scala 29:58]
  assign _T_2085 = _T_2059[3:0]; // @[LZD.scala 44:32]
  assign _T_2086 = _T_2085[3:2]; // @[LZD.scala 43:32]
  assign _T_2087 = _T_2086 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2088 = _T_2086[1]; // @[LZD.scala 39:21]
  assign _T_2089 = _T_2086[0]; // @[LZD.scala 39:30]
  assign _T_2090 = ~ _T_2089; // @[LZD.scala 39:27]
  assign _T_2091 = _T_2088 | _T_2090; // @[LZD.scala 39:25]
  assign _T_2092 = {_T_2087,_T_2091}; // @[Cat.scala 29:58]
  assign _T_2093 = _T_2085[1:0]; // @[LZD.scala 44:32]
  assign _T_2094 = _T_2093 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2095 = _T_2093[1]; // @[LZD.scala 39:21]
  assign _T_2096 = _T_2093[0]; // @[LZD.scala 39:30]
  assign _T_2097 = ~ _T_2096; // @[LZD.scala 39:27]
  assign _T_2098 = _T_2095 | _T_2097; // @[LZD.scala 39:25]
  assign _T_2099 = {_T_2094,_T_2098}; // @[Cat.scala 29:58]
  assign _T_2100 = _T_2092[1]; // @[Shift.scala 12:21]
  assign _T_2101 = _T_2099[1]; // @[Shift.scala 12:21]
  assign _T_2102 = _T_2100 | _T_2101; // @[LZD.scala 49:16]
  assign _T_2103 = ~ _T_2101; // @[LZD.scala 49:27]
  assign _T_2104 = _T_2100 | _T_2103; // @[LZD.scala 49:25]
  assign _T_2105 = _T_2092[0:0]; // @[LZD.scala 49:47]
  assign _T_2106 = _T_2099[0:0]; // @[LZD.scala 49:59]
  assign _T_2107 = _T_2100 ? _T_2105 : _T_2106; // @[LZD.scala 49:35]
  assign _T_2109 = {_T_2102,_T_2104,_T_2107}; // @[Cat.scala 29:58]
  assign _T_2110 = _T_2084[2]; // @[Shift.scala 12:21]
  assign _T_2111 = _T_2109[2]; // @[Shift.scala 12:21]
  assign _T_2112 = _T_2110 | _T_2111; // @[LZD.scala 49:16]
  assign _T_2113 = ~ _T_2111; // @[LZD.scala 49:27]
  assign _T_2114 = _T_2110 | _T_2113; // @[LZD.scala 49:25]
  assign _T_2115 = _T_2084[1:0]; // @[LZD.scala 49:47]
  assign _T_2116 = _T_2109[1:0]; // @[LZD.scala 49:59]
  assign _T_2117 = _T_2110 ? _T_2115 : _T_2116; // @[LZD.scala 49:35]
  assign _T_2119 = {_T_2112,_T_2114,_T_2117}; // @[Cat.scala 29:58]
  assign _T_2120 = _T_2058[3]; // @[Shift.scala 12:21]
  assign _T_2121 = _T_2119[3]; // @[Shift.scala 12:21]
  assign _T_2122 = _T_2120 | _T_2121; // @[LZD.scala 49:16]
  assign _T_2123 = ~ _T_2121; // @[LZD.scala 49:27]
  assign _T_2124 = _T_2120 | _T_2123; // @[LZD.scala 49:25]
  assign _T_2125 = _T_2058[2:0]; // @[LZD.scala 49:47]
  assign _T_2126 = _T_2119[2:0]; // @[LZD.scala 49:59]
  assign _T_2127 = _T_2120 ? _T_2125 : _T_2126; // @[LZD.scala 49:35]
  assign _T_2129 = {_T_2122,_T_2124,_T_2127}; // @[Cat.scala 29:58]
  assign _T_2130 = _T_1996[15:0]; // @[LZD.scala 44:32]
  assign _T_2131 = _T_2130[15:8]; // @[LZD.scala 43:32]
  assign _T_2132 = _T_2131[7:4]; // @[LZD.scala 43:32]
  assign _T_2133 = _T_2132[3:2]; // @[LZD.scala 43:32]
  assign _T_2134 = _T_2133 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2135 = _T_2133[1]; // @[LZD.scala 39:21]
  assign _T_2136 = _T_2133[0]; // @[LZD.scala 39:30]
  assign _T_2137 = ~ _T_2136; // @[LZD.scala 39:27]
  assign _T_2138 = _T_2135 | _T_2137; // @[LZD.scala 39:25]
  assign _T_2139 = {_T_2134,_T_2138}; // @[Cat.scala 29:58]
  assign _T_2140 = _T_2132[1:0]; // @[LZD.scala 44:32]
  assign _T_2141 = _T_2140 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2142 = _T_2140[1]; // @[LZD.scala 39:21]
  assign _T_2143 = _T_2140[0]; // @[LZD.scala 39:30]
  assign _T_2144 = ~ _T_2143; // @[LZD.scala 39:27]
  assign _T_2145 = _T_2142 | _T_2144; // @[LZD.scala 39:25]
  assign _T_2146 = {_T_2141,_T_2145}; // @[Cat.scala 29:58]
  assign _T_2147 = _T_2139[1]; // @[Shift.scala 12:21]
  assign _T_2148 = _T_2146[1]; // @[Shift.scala 12:21]
  assign _T_2149 = _T_2147 | _T_2148; // @[LZD.scala 49:16]
  assign _T_2150 = ~ _T_2148; // @[LZD.scala 49:27]
  assign _T_2151 = _T_2147 | _T_2150; // @[LZD.scala 49:25]
  assign _T_2152 = _T_2139[0:0]; // @[LZD.scala 49:47]
  assign _T_2153 = _T_2146[0:0]; // @[LZD.scala 49:59]
  assign _T_2154 = _T_2147 ? _T_2152 : _T_2153; // @[LZD.scala 49:35]
  assign _T_2156 = {_T_2149,_T_2151,_T_2154}; // @[Cat.scala 29:58]
  assign _T_2157 = _T_2131[3:0]; // @[LZD.scala 44:32]
  assign _T_2158 = _T_2157[3:2]; // @[LZD.scala 43:32]
  assign _T_2159 = _T_2158 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2160 = _T_2158[1]; // @[LZD.scala 39:21]
  assign _T_2161 = _T_2158[0]; // @[LZD.scala 39:30]
  assign _T_2162 = ~ _T_2161; // @[LZD.scala 39:27]
  assign _T_2163 = _T_2160 | _T_2162; // @[LZD.scala 39:25]
  assign _T_2164 = {_T_2159,_T_2163}; // @[Cat.scala 29:58]
  assign _T_2165 = _T_2157[1:0]; // @[LZD.scala 44:32]
  assign _T_2166 = _T_2165 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2167 = _T_2165[1]; // @[LZD.scala 39:21]
  assign _T_2168 = _T_2165[0]; // @[LZD.scala 39:30]
  assign _T_2169 = ~ _T_2168; // @[LZD.scala 39:27]
  assign _T_2170 = _T_2167 | _T_2169; // @[LZD.scala 39:25]
  assign _T_2171 = {_T_2166,_T_2170}; // @[Cat.scala 29:58]
  assign _T_2172 = _T_2164[1]; // @[Shift.scala 12:21]
  assign _T_2173 = _T_2171[1]; // @[Shift.scala 12:21]
  assign _T_2174 = _T_2172 | _T_2173; // @[LZD.scala 49:16]
  assign _T_2175 = ~ _T_2173; // @[LZD.scala 49:27]
  assign _T_2176 = _T_2172 | _T_2175; // @[LZD.scala 49:25]
  assign _T_2177 = _T_2164[0:0]; // @[LZD.scala 49:47]
  assign _T_2178 = _T_2171[0:0]; // @[LZD.scala 49:59]
  assign _T_2179 = _T_2172 ? _T_2177 : _T_2178; // @[LZD.scala 49:35]
  assign _T_2181 = {_T_2174,_T_2176,_T_2179}; // @[Cat.scala 29:58]
  assign _T_2182 = _T_2156[2]; // @[Shift.scala 12:21]
  assign _T_2183 = _T_2181[2]; // @[Shift.scala 12:21]
  assign _T_2184 = _T_2182 | _T_2183; // @[LZD.scala 49:16]
  assign _T_2185 = ~ _T_2183; // @[LZD.scala 49:27]
  assign _T_2186 = _T_2182 | _T_2185; // @[LZD.scala 49:25]
  assign _T_2187 = _T_2156[1:0]; // @[LZD.scala 49:47]
  assign _T_2188 = _T_2181[1:0]; // @[LZD.scala 49:59]
  assign _T_2189 = _T_2182 ? _T_2187 : _T_2188; // @[LZD.scala 49:35]
  assign _T_2191 = {_T_2184,_T_2186,_T_2189}; // @[Cat.scala 29:58]
  assign _T_2192 = _T_2130[7:0]; // @[LZD.scala 44:32]
  assign _T_2193 = _T_2192[7:4]; // @[LZD.scala 43:32]
  assign _T_2194 = _T_2193[3:2]; // @[LZD.scala 43:32]
  assign _T_2195 = _T_2194 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2196 = _T_2194[1]; // @[LZD.scala 39:21]
  assign _T_2197 = _T_2194[0]; // @[LZD.scala 39:30]
  assign _T_2198 = ~ _T_2197; // @[LZD.scala 39:27]
  assign _T_2199 = _T_2196 | _T_2198; // @[LZD.scala 39:25]
  assign _T_2200 = {_T_2195,_T_2199}; // @[Cat.scala 29:58]
  assign _T_2201 = _T_2193[1:0]; // @[LZD.scala 44:32]
  assign _T_2202 = _T_2201 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2203 = _T_2201[1]; // @[LZD.scala 39:21]
  assign _T_2204 = _T_2201[0]; // @[LZD.scala 39:30]
  assign _T_2205 = ~ _T_2204; // @[LZD.scala 39:27]
  assign _T_2206 = _T_2203 | _T_2205; // @[LZD.scala 39:25]
  assign _T_2207 = {_T_2202,_T_2206}; // @[Cat.scala 29:58]
  assign _T_2208 = _T_2200[1]; // @[Shift.scala 12:21]
  assign _T_2209 = _T_2207[1]; // @[Shift.scala 12:21]
  assign _T_2210 = _T_2208 | _T_2209; // @[LZD.scala 49:16]
  assign _T_2211 = ~ _T_2209; // @[LZD.scala 49:27]
  assign _T_2212 = _T_2208 | _T_2211; // @[LZD.scala 49:25]
  assign _T_2213 = _T_2200[0:0]; // @[LZD.scala 49:47]
  assign _T_2214 = _T_2207[0:0]; // @[LZD.scala 49:59]
  assign _T_2215 = _T_2208 ? _T_2213 : _T_2214; // @[LZD.scala 49:35]
  assign _T_2217 = {_T_2210,_T_2212,_T_2215}; // @[Cat.scala 29:58]
  assign _T_2218 = _T_2192[3:0]; // @[LZD.scala 44:32]
  assign _T_2219 = _T_2218[3:2]; // @[LZD.scala 43:32]
  assign _T_2220 = _T_2219 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2221 = _T_2219[1]; // @[LZD.scala 39:21]
  assign _T_2222 = _T_2219[0]; // @[LZD.scala 39:30]
  assign _T_2223 = ~ _T_2222; // @[LZD.scala 39:27]
  assign _T_2224 = _T_2221 | _T_2223; // @[LZD.scala 39:25]
  assign _T_2225 = {_T_2220,_T_2224}; // @[Cat.scala 29:58]
  assign _T_2226 = _T_2218[1:0]; // @[LZD.scala 44:32]
  assign _T_2227 = _T_2226 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2228 = _T_2226[1]; // @[LZD.scala 39:21]
  assign _T_2229 = _T_2226[0]; // @[LZD.scala 39:30]
  assign _T_2230 = ~ _T_2229; // @[LZD.scala 39:27]
  assign _T_2231 = _T_2228 | _T_2230; // @[LZD.scala 39:25]
  assign _T_2232 = {_T_2227,_T_2231}; // @[Cat.scala 29:58]
  assign _T_2233 = _T_2225[1]; // @[Shift.scala 12:21]
  assign _T_2234 = _T_2232[1]; // @[Shift.scala 12:21]
  assign _T_2235 = _T_2233 | _T_2234; // @[LZD.scala 49:16]
  assign _T_2236 = ~ _T_2234; // @[LZD.scala 49:27]
  assign _T_2237 = _T_2233 | _T_2236; // @[LZD.scala 49:25]
  assign _T_2238 = _T_2225[0:0]; // @[LZD.scala 49:47]
  assign _T_2239 = _T_2232[0:0]; // @[LZD.scala 49:59]
  assign _T_2240 = _T_2233 ? _T_2238 : _T_2239; // @[LZD.scala 49:35]
  assign _T_2242 = {_T_2235,_T_2237,_T_2240}; // @[Cat.scala 29:58]
  assign _T_2243 = _T_2217[2]; // @[Shift.scala 12:21]
  assign _T_2244 = _T_2242[2]; // @[Shift.scala 12:21]
  assign _T_2245 = _T_2243 | _T_2244; // @[LZD.scala 49:16]
  assign _T_2246 = ~ _T_2244; // @[LZD.scala 49:27]
  assign _T_2247 = _T_2243 | _T_2246; // @[LZD.scala 49:25]
  assign _T_2248 = _T_2217[1:0]; // @[LZD.scala 49:47]
  assign _T_2249 = _T_2242[1:0]; // @[LZD.scala 49:59]
  assign _T_2250 = _T_2243 ? _T_2248 : _T_2249; // @[LZD.scala 49:35]
  assign _T_2252 = {_T_2245,_T_2247,_T_2250}; // @[Cat.scala 29:58]
  assign _T_2253 = _T_2191[3]; // @[Shift.scala 12:21]
  assign _T_2254 = _T_2252[3]; // @[Shift.scala 12:21]
  assign _T_2255 = _T_2253 | _T_2254; // @[LZD.scala 49:16]
  assign _T_2256 = ~ _T_2254; // @[LZD.scala 49:27]
  assign _T_2257 = _T_2253 | _T_2256; // @[LZD.scala 49:25]
  assign _T_2258 = _T_2191[2:0]; // @[LZD.scala 49:47]
  assign _T_2259 = _T_2252[2:0]; // @[LZD.scala 49:59]
  assign _T_2260 = _T_2253 ? _T_2258 : _T_2259; // @[LZD.scala 49:35]
  assign _T_2262 = {_T_2255,_T_2257,_T_2260}; // @[Cat.scala 29:58]
  assign _T_2263 = _T_2129[4]; // @[Shift.scala 12:21]
  assign _T_2264 = _T_2262[4]; // @[Shift.scala 12:21]
  assign _T_2265 = _T_2263 | _T_2264; // @[LZD.scala 49:16]
  assign _T_2266 = ~ _T_2264; // @[LZD.scala 49:27]
  assign _T_2267 = _T_2263 | _T_2266; // @[LZD.scala 49:25]
  assign _T_2268 = _T_2129[3:0]; // @[LZD.scala 49:47]
  assign _T_2269 = _T_2262[3:0]; // @[LZD.scala 49:59]
  assign _T_2270 = _T_2263 ? _T_2268 : _T_2269; // @[LZD.scala 49:35]
  assign _T_2272 = {_T_2265,_T_2267,_T_2270}; // @[Cat.scala 29:58]
  assign _T_2273 = _T_1995[5]; // @[Shift.scala 12:21]
  assign _T_2274 = _T_2272[5]; // @[Shift.scala 12:21]
  assign _T_2275 = _T_2273 | _T_2274; // @[LZD.scala 49:16]
  assign _T_2276 = ~ _T_2274; // @[LZD.scala 49:27]
  assign _T_2277 = _T_2273 | _T_2276; // @[LZD.scala 49:25]
  assign _T_2278 = _T_1995[4:0]; // @[LZD.scala 49:47]
  assign _T_2279 = _T_2272[4:0]; // @[LZD.scala 49:59]
  assign _T_2280 = _T_2273 ? _T_2278 : _T_2279; // @[LZD.scala 49:35]
  assign _T_2282 = {_T_2275,_T_2277,_T_2280}; // @[Cat.scala 29:58]
  assign _T_2283 = _T_1717[6]; // @[Shift.scala 12:21]
  assign _T_2284 = _T_2282[6]; // @[Shift.scala 12:21]
  assign _T_2285 = _T_2283 | _T_2284; // @[LZD.scala 49:16]
  assign _T_2286 = ~ _T_2284; // @[LZD.scala 49:27]
  assign _T_2287 = _T_2283 | _T_2286; // @[LZD.scala 49:25]
  assign _T_2288 = _T_1717[5:0]; // @[LZD.scala 49:47]
  assign _T_2289 = _T_2282[5:0]; // @[LZD.scala 49:59]
  assign _T_2290 = _T_2283 ? _T_2288 : _T_2289; // @[LZD.scala 49:35]
  assign _T_2292 = {_T_2285,_T_2287,_T_2290}; // @[Cat.scala 29:58]
  assign _T_2293 = _T_1151[7]; // @[Shift.scala 12:21]
  assign _T_2294 = _T_2292[7]; // @[Shift.scala 12:21]
  assign _T_2295 = _T_2293 | _T_2294; // @[LZD.scala 49:16]
  assign _T_2296 = ~ _T_2294; // @[LZD.scala 49:27]
  assign _T_2297 = _T_2293 | _T_2296; // @[LZD.scala 49:25]
  assign _T_2298 = _T_1151[6:0]; // @[LZD.scala 49:47]
  assign _T_2299 = _T_2292[6:0]; // @[LZD.scala 49:59]
  assign _T_2300 = _T_2293 ? _T_2298 : _T_2299; // @[LZD.scala 49:35]
  assign _T_2302 = {_T_2295,_T_2297,_T_2300}; // @[Cat.scala 29:58]
  assign _T_2303 = quireXOR[56:0]; // @[LZD.scala 44:32]
  assign _T_2304 = _T_2303[56:25]; // @[LZD.scala 43:32]
  assign _T_2305 = _T_2304[31:16]; // @[LZD.scala 43:32]
  assign _T_2306 = _T_2305[15:8]; // @[LZD.scala 43:32]
  assign _T_2307 = _T_2306[7:4]; // @[LZD.scala 43:32]
  assign _T_2308 = _T_2307[3:2]; // @[LZD.scala 43:32]
  assign _T_2309 = _T_2308 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2310 = _T_2308[1]; // @[LZD.scala 39:21]
  assign _T_2311 = _T_2308[0]; // @[LZD.scala 39:30]
  assign _T_2312 = ~ _T_2311; // @[LZD.scala 39:27]
  assign _T_2313 = _T_2310 | _T_2312; // @[LZD.scala 39:25]
  assign _T_2314 = {_T_2309,_T_2313}; // @[Cat.scala 29:58]
  assign _T_2315 = _T_2307[1:0]; // @[LZD.scala 44:32]
  assign _T_2316 = _T_2315 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2317 = _T_2315[1]; // @[LZD.scala 39:21]
  assign _T_2318 = _T_2315[0]; // @[LZD.scala 39:30]
  assign _T_2319 = ~ _T_2318; // @[LZD.scala 39:27]
  assign _T_2320 = _T_2317 | _T_2319; // @[LZD.scala 39:25]
  assign _T_2321 = {_T_2316,_T_2320}; // @[Cat.scala 29:58]
  assign _T_2322 = _T_2314[1]; // @[Shift.scala 12:21]
  assign _T_2323 = _T_2321[1]; // @[Shift.scala 12:21]
  assign _T_2324 = _T_2322 | _T_2323; // @[LZD.scala 49:16]
  assign _T_2325 = ~ _T_2323; // @[LZD.scala 49:27]
  assign _T_2326 = _T_2322 | _T_2325; // @[LZD.scala 49:25]
  assign _T_2327 = _T_2314[0:0]; // @[LZD.scala 49:47]
  assign _T_2328 = _T_2321[0:0]; // @[LZD.scala 49:59]
  assign _T_2329 = _T_2322 ? _T_2327 : _T_2328; // @[LZD.scala 49:35]
  assign _T_2331 = {_T_2324,_T_2326,_T_2329}; // @[Cat.scala 29:58]
  assign _T_2332 = _T_2306[3:0]; // @[LZD.scala 44:32]
  assign _T_2333 = _T_2332[3:2]; // @[LZD.scala 43:32]
  assign _T_2334 = _T_2333 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2335 = _T_2333[1]; // @[LZD.scala 39:21]
  assign _T_2336 = _T_2333[0]; // @[LZD.scala 39:30]
  assign _T_2337 = ~ _T_2336; // @[LZD.scala 39:27]
  assign _T_2338 = _T_2335 | _T_2337; // @[LZD.scala 39:25]
  assign _T_2339 = {_T_2334,_T_2338}; // @[Cat.scala 29:58]
  assign _T_2340 = _T_2332[1:0]; // @[LZD.scala 44:32]
  assign _T_2341 = _T_2340 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2342 = _T_2340[1]; // @[LZD.scala 39:21]
  assign _T_2343 = _T_2340[0]; // @[LZD.scala 39:30]
  assign _T_2344 = ~ _T_2343; // @[LZD.scala 39:27]
  assign _T_2345 = _T_2342 | _T_2344; // @[LZD.scala 39:25]
  assign _T_2346 = {_T_2341,_T_2345}; // @[Cat.scala 29:58]
  assign _T_2347 = _T_2339[1]; // @[Shift.scala 12:21]
  assign _T_2348 = _T_2346[1]; // @[Shift.scala 12:21]
  assign _T_2349 = _T_2347 | _T_2348; // @[LZD.scala 49:16]
  assign _T_2350 = ~ _T_2348; // @[LZD.scala 49:27]
  assign _T_2351 = _T_2347 | _T_2350; // @[LZD.scala 49:25]
  assign _T_2352 = _T_2339[0:0]; // @[LZD.scala 49:47]
  assign _T_2353 = _T_2346[0:0]; // @[LZD.scala 49:59]
  assign _T_2354 = _T_2347 ? _T_2352 : _T_2353; // @[LZD.scala 49:35]
  assign _T_2356 = {_T_2349,_T_2351,_T_2354}; // @[Cat.scala 29:58]
  assign _T_2357 = _T_2331[2]; // @[Shift.scala 12:21]
  assign _T_2358 = _T_2356[2]; // @[Shift.scala 12:21]
  assign _T_2359 = _T_2357 | _T_2358; // @[LZD.scala 49:16]
  assign _T_2360 = ~ _T_2358; // @[LZD.scala 49:27]
  assign _T_2361 = _T_2357 | _T_2360; // @[LZD.scala 49:25]
  assign _T_2362 = _T_2331[1:0]; // @[LZD.scala 49:47]
  assign _T_2363 = _T_2356[1:0]; // @[LZD.scala 49:59]
  assign _T_2364 = _T_2357 ? _T_2362 : _T_2363; // @[LZD.scala 49:35]
  assign _T_2366 = {_T_2359,_T_2361,_T_2364}; // @[Cat.scala 29:58]
  assign _T_2367 = _T_2305[7:0]; // @[LZD.scala 44:32]
  assign _T_2368 = _T_2367[7:4]; // @[LZD.scala 43:32]
  assign _T_2369 = _T_2368[3:2]; // @[LZD.scala 43:32]
  assign _T_2370 = _T_2369 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2371 = _T_2369[1]; // @[LZD.scala 39:21]
  assign _T_2372 = _T_2369[0]; // @[LZD.scala 39:30]
  assign _T_2373 = ~ _T_2372; // @[LZD.scala 39:27]
  assign _T_2374 = _T_2371 | _T_2373; // @[LZD.scala 39:25]
  assign _T_2375 = {_T_2370,_T_2374}; // @[Cat.scala 29:58]
  assign _T_2376 = _T_2368[1:0]; // @[LZD.scala 44:32]
  assign _T_2377 = _T_2376 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2378 = _T_2376[1]; // @[LZD.scala 39:21]
  assign _T_2379 = _T_2376[0]; // @[LZD.scala 39:30]
  assign _T_2380 = ~ _T_2379; // @[LZD.scala 39:27]
  assign _T_2381 = _T_2378 | _T_2380; // @[LZD.scala 39:25]
  assign _T_2382 = {_T_2377,_T_2381}; // @[Cat.scala 29:58]
  assign _T_2383 = _T_2375[1]; // @[Shift.scala 12:21]
  assign _T_2384 = _T_2382[1]; // @[Shift.scala 12:21]
  assign _T_2385 = _T_2383 | _T_2384; // @[LZD.scala 49:16]
  assign _T_2386 = ~ _T_2384; // @[LZD.scala 49:27]
  assign _T_2387 = _T_2383 | _T_2386; // @[LZD.scala 49:25]
  assign _T_2388 = _T_2375[0:0]; // @[LZD.scala 49:47]
  assign _T_2389 = _T_2382[0:0]; // @[LZD.scala 49:59]
  assign _T_2390 = _T_2383 ? _T_2388 : _T_2389; // @[LZD.scala 49:35]
  assign _T_2392 = {_T_2385,_T_2387,_T_2390}; // @[Cat.scala 29:58]
  assign _T_2393 = _T_2367[3:0]; // @[LZD.scala 44:32]
  assign _T_2394 = _T_2393[3:2]; // @[LZD.scala 43:32]
  assign _T_2395 = _T_2394 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2396 = _T_2394[1]; // @[LZD.scala 39:21]
  assign _T_2397 = _T_2394[0]; // @[LZD.scala 39:30]
  assign _T_2398 = ~ _T_2397; // @[LZD.scala 39:27]
  assign _T_2399 = _T_2396 | _T_2398; // @[LZD.scala 39:25]
  assign _T_2400 = {_T_2395,_T_2399}; // @[Cat.scala 29:58]
  assign _T_2401 = _T_2393[1:0]; // @[LZD.scala 44:32]
  assign _T_2402 = _T_2401 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2403 = _T_2401[1]; // @[LZD.scala 39:21]
  assign _T_2404 = _T_2401[0]; // @[LZD.scala 39:30]
  assign _T_2405 = ~ _T_2404; // @[LZD.scala 39:27]
  assign _T_2406 = _T_2403 | _T_2405; // @[LZD.scala 39:25]
  assign _T_2407 = {_T_2402,_T_2406}; // @[Cat.scala 29:58]
  assign _T_2408 = _T_2400[1]; // @[Shift.scala 12:21]
  assign _T_2409 = _T_2407[1]; // @[Shift.scala 12:21]
  assign _T_2410 = _T_2408 | _T_2409; // @[LZD.scala 49:16]
  assign _T_2411 = ~ _T_2409; // @[LZD.scala 49:27]
  assign _T_2412 = _T_2408 | _T_2411; // @[LZD.scala 49:25]
  assign _T_2413 = _T_2400[0:0]; // @[LZD.scala 49:47]
  assign _T_2414 = _T_2407[0:0]; // @[LZD.scala 49:59]
  assign _T_2415 = _T_2408 ? _T_2413 : _T_2414; // @[LZD.scala 49:35]
  assign _T_2417 = {_T_2410,_T_2412,_T_2415}; // @[Cat.scala 29:58]
  assign _T_2418 = _T_2392[2]; // @[Shift.scala 12:21]
  assign _T_2419 = _T_2417[2]; // @[Shift.scala 12:21]
  assign _T_2420 = _T_2418 | _T_2419; // @[LZD.scala 49:16]
  assign _T_2421 = ~ _T_2419; // @[LZD.scala 49:27]
  assign _T_2422 = _T_2418 | _T_2421; // @[LZD.scala 49:25]
  assign _T_2423 = _T_2392[1:0]; // @[LZD.scala 49:47]
  assign _T_2424 = _T_2417[1:0]; // @[LZD.scala 49:59]
  assign _T_2425 = _T_2418 ? _T_2423 : _T_2424; // @[LZD.scala 49:35]
  assign _T_2427 = {_T_2420,_T_2422,_T_2425}; // @[Cat.scala 29:58]
  assign _T_2428 = _T_2366[3]; // @[Shift.scala 12:21]
  assign _T_2429 = _T_2427[3]; // @[Shift.scala 12:21]
  assign _T_2430 = _T_2428 | _T_2429; // @[LZD.scala 49:16]
  assign _T_2431 = ~ _T_2429; // @[LZD.scala 49:27]
  assign _T_2432 = _T_2428 | _T_2431; // @[LZD.scala 49:25]
  assign _T_2433 = _T_2366[2:0]; // @[LZD.scala 49:47]
  assign _T_2434 = _T_2427[2:0]; // @[LZD.scala 49:59]
  assign _T_2435 = _T_2428 ? _T_2433 : _T_2434; // @[LZD.scala 49:35]
  assign _T_2437 = {_T_2430,_T_2432,_T_2435}; // @[Cat.scala 29:58]
  assign _T_2438 = _T_2304[15:0]; // @[LZD.scala 44:32]
  assign _T_2439 = _T_2438[15:8]; // @[LZD.scala 43:32]
  assign _T_2440 = _T_2439[7:4]; // @[LZD.scala 43:32]
  assign _T_2441 = _T_2440[3:2]; // @[LZD.scala 43:32]
  assign _T_2442 = _T_2441 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2443 = _T_2441[1]; // @[LZD.scala 39:21]
  assign _T_2444 = _T_2441[0]; // @[LZD.scala 39:30]
  assign _T_2445 = ~ _T_2444; // @[LZD.scala 39:27]
  assign _T_2446 = _T_2443 | _T_2445; // @[LZD.scala 39:25]
  assign _T_2447 = {_T_2442,_T_2446}; // @[Cat.scala 29:58]
  assign _T_2448 = _T_2440[1:0]; // @[LZD.scala 44:32]
  assign _T_2449 = _T_2448 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2450 = _T_2448[1]; // @[LZD.scala 39:21]
  assign _T_2451 = _T_2448[0]; // @[LZD.scala 39:30]
  assign _T_2452 = ~ _T_2451; // @[LZD.scala 39:27]
  assign _T_2453 = _T_2450 | _T_2452; // @[LZD.scala 39:25]
  assign _T_2454 = {_T_2449,_T_2453}; // @[Cat.scala 29:58]
  assign _T_2455 = _T_2447[1]; // @[Shift.scala 12:21]
  assign _T_2456 = _T_2454[1]; // @[Shift.scala 12:21]
  assign _T_2457 = _T_2455 | _T_2456; // @[LZD.scala 49:16]
  assign _T_2458 = ~ _T_2456; // @[LZD.scala 49:27]
  assign _T_2459 = _T_2455 | _T_2458; // @[LZD.scala 49:25]
  assign _T_2460 = _T_2447[0:0]; // @[LZD.scala 49:47]
  assign _T_2461 = _T_2454[0:0]; // @[LZD.scala 49:59]
  assign _T_2462 = _T_2455 ? _T_2460 : _T_2461; // @[LZD.scala 49:35]
  assign _T_2464 = {_T_2457,_T_2459,_T_2462}; // @[Cat.scala 29:58]
  assign _T_2465 = _T_2439[3:0]; // @[LZD.scala 44:32]
  assign _T_2466 = _T_2465[3:2]; // @[LZD.scala 43:32]
  assign _T_2467 = _T_2466 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2468 = _T_2466[1]; // @[LZD.scala 39:21]
  assign _T_2469 = _T_2466[0]; // @[LZD.scala 39:30]
  assign _T_2470 = ~ _T_2469; // @[LZD.scala 39:27]
  assign _T_2471 = _T_2468 | _T_2470; // @[LZD.scala 39:25]
  assign _T_2472 = {_T_2467,_T_2471}; // @[Cat.scala 29:58]
  assign _T_2473 = _T_2465[1:0]; // @[LZD.scala 44:32]
  assign _T_2474 = _T_2473 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2475 = _T_2473[1]; // @[LZD.scala 39:21]
  assign _T_2476 = _T_2473[0]; // @[LZD.scala 39:30]
  assign _T_2477 = ~ _T_2476; // @[LZD.scala 39:27]
  assign _T_2478 = _T_2475 | _T_2477; // @[LZD.scala 39:25]
  assign _T_2479 = {_T_2474,_T_2478}; // @[Cat.scala 29:58]
  assign _T_2480 = _T_2472[1]; // @[Shift.scala 12:21]
  assign _T_2481 = _T_2479[1]; // @[Shift.scala 12:21]
  assign _T_2482 = _T_2480 | _T_2481; // @[LZD.scala 49:16]
  assign _T_2483 = ~ _T_2481; // @[LZD.scala 49:27]
  assign _T_2484 = _T_2480 | _T_2483; // @[LZD.scala 49:25]
  assign _T_2485 = _T_2472[0:0]; // @[LZD.scala 49:47]
  assign _T_2486 = _T_2479[0:0]; // @[LZD.scala 49:59]
  assign _T_2487 = _T_2480 ? _T_2485 : _T_2486; // @[LZD.scala 49:35]
  assign _T_2489 = {_T_2482,_T_2484,_T_2487}; // @[Cat.scala 29:58]
  assign _T_2490 = _T_2464[2]; // @[Shift.scala 12:21]
  assign _T_2491 = _T_2489[2]; // @[Shift.scala 12:21]
  assign _T_2492 = _T_2490 | _T_2491; // @[LZD.scala 49:16]
  assign _T_2493 = ~ _T_2491; // @[LZD.scala 49:27]
  assign _T_2494 = _T_2490 | _T_2493; // @[LZD.scala 49:25]
  assign _T_2495 = _T_2464[1:0]; // @[LZD.scala 49:47]
  assign _T_2496 = _T_2489[1:0]; // @[LZD.scala 49:59]
  assign _T_2497 = _T_2490 ? _T_2495 : _T_2496; // @[LZD.scala 49:35]
  assign _T_2499 = {_T_2492,_T_2494,_T_2497}; // @[Cat.scala 29:58]
  assign _T_2500 = _T_2438[7:0]; // @[LZD.scala 44:32]
  assign _T_2501 = _T_2500[7:4]; // @[LZD.scala 43:32]
  assign _T_2502 = _T_2501[3:2]; // @[LZD.scala 43:32]
  assign _T_2503 = _T_2502 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2504 = _T_2502[1]; // @[LZD.scala 39:21]
  assign _T_2505 = _T_2502[0]; // @[LZD.scala 39:30]
  assign _T_2506 = ~ _T_2505; // @[LZD.scala 39:27]
  assign _T_2507 = _T_2504 | _T_2506; // @[LZD.scala 39:25]
  assign _T_2508 = {_T_2503,_T_2507}; // @[Cat.scala 29:58]
  assign _T_2509 = _T_2501[1:0]; // @[LZD.scala 44:32]
  assign _T_2510 = _T_2509 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2511 = _T_2509[1]; // @[LZD.scala 39:21]
  assign _T_2512 = _T_2509[0]; // @[LZD.scala 39:30]
  assign _T_2513 = ~ _T_2512; // @[LZD.scala 39:27]
  assign _T_2514 = _T_2511 | _T_2513; // @[LZD.scala 39:25]
  assign _T_2515 = {_T_2510,_T_2514}; // @[Cat.scala 29:58]
  assign _T_2516 = _T_2508[1]; // @[Shift.scala 12:21]
  assign _T_2517 = _T_2515[1]; // @[Shift.scala 12:21]
  assign _T_2518 = _T_2516 | _T_2517; // @[LZD.scala 49:16]
  assign _T_2519 = ~ _T_2517; // @[LZD.scala 49:27]
  assign _T_2520 = _T_2516 | _T_2519; // @[LZD.scala 49:25]
  assign _T_2521 = _T_2508[0:0]; // @[LZD.scala 49:47]
  assign _T_2522 = _T_2515[0:0]; // @[LZD.scala 49:59]
  assign _T_2523 = _T_2516 ? _T_2521 : _T_2522; // @[LZD.scala 49:35]
  assign _T_2525 = {_T_2518,_T_2520,_T_2523}; // @[Cat.scala 29:58]
  assign _T_2526 = _T_2500[3:0]; // @[LZD.scala 44:32]
  assign _T_2527 = _T_2526[3:2]; // @[LZD.scala 43:32]
  assign _T_2528 = _T_2527 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2529 = _T_2527[1]; // @[LZD.scala 39:21]
  assign _T_2530 = _T_2527[0]; // @[LZD.scala 39:30]
  assign _T_2531 = ~ _T_2530; // @[LZD.scala 39:27]
  assign _T_2532 = _T_2529 | _T_2531; // @[LZD.scala 39:25]
  assign _T_2533 = {_T_2528,_T_2532}; // @[Cat.scala 29:58]
  assign _T_2534 = _T_2526[1:0]; // @[LZD.scala 44:32]
  assign _T_2535 = _T_2534 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2536 = _T_2534[1]; // @[LZD.scala 39:21]
  assign _T_2537 = _T_2534[0]; // @[LZD.scala 39:30]
  assign _T_2538 = ~ _T_2537; // @[LZD.scala 39:27]
  assign _T_2539 = _T_2536 | _T_2538; // @[LZD.scala 39:25]
  assign _T_2540 = {_T_2535,_T_2539}; // @[Cat.scala 29:58]
  assign _T_2541 = _T_2533[1]; // @[Shift.scala 12:21]
  assign _T_2542 = _T_2540[1]; // @[Shift.scala 12:21]
  assign _T_2543 = _T_2541 | _T_2542; // @[LZD.scala 49:16]
  assign _T_2544 = ~ _T_2542; // @[LZD.scala 49:27]
  assign _T_2545 = _T_2541 | _T_2544; // @[LZD.scala 49:25]
  assign _T_2546 = _T_2533[0:0]; // @[LZD.scala 49:47]
  assign _T_2547 = _T_2540[0:0]; // @[LZD.scala 49:59]
  assign _T_2548 = _T_2541 ? _T_2546 : _T_2547; // @[LZD.scala 49:35]
  assign _T_2550 = {_T_2543,_T_2545,_T_2548}; // @[Cat.scala 29:58]
  assign _T_2551 = _T_2525[2]; // @[Shift.scala 12:21]
  assign _T_2552 = _T_2550[2]; // @[Shift.scala 12:21]
  assign _T_2553 = _T_2551 | _T_2552; // @[LZD.scala 49:16]
  assign _T_2554 = ~ _T_2552; // @[LZD.scala 49:27]
  assign _T_2555 = _T_2551 | _T_2554; // @[LZD.scala 49:25]
  assign _T_2556 = _T_2525[1:0]; // @[LZD.scala 49:47]
  assign _T_2557 = _T_2550[1:0]; // @[LZD.scala 49:59]
  assign _T_2558 = _T_2551 ? _T_2556 : _T_2557; // @[LZD.scala 49:35]
  assign _T_2560 = {_T_2553,_T_2555,_T_2558}; // @[Cat.scala 29:58]
  assign _T_2561 = _T_2499[3]; // @[Shift.scala 12:21]
  assign _T_2562 = _T_2560[3]; // @[Shift.scala 12:21]
  assign _T_2563 = _T_2561 | _T_2562; // @[LZD.scala 49:16]
  assign _T_2564 = ~ _T_2562; // @[LZD.scala 49:27]
  assign _T_2565 = _T_2561 | _T_2564; // @[LZD.scala 49:25]
  assign _T_2566 = _T_2499[2:0]; // @[LZD.scala 49:47]
  assign _T_2567 = _T_2560[2:0]; // @[LZD.scala 49:59]
  assign _T_2568 = _T_2561 ? _T_2566 : _T_2567; // @[LZD.scala 49:35]
  assign _T_2570 = {_T_2563,_T_2565,_T_2568}; // @[Cat.scala 29:58]
  assign _T_2571 = _T_2437[4]; // @[Shift.scala 12:21]
  assign _T_2572 = _T_2570[4]; // @[Shift.scala 12:21]
  assign _T_2573 = _T_2571 | _T_2572; // @[LZD.scala 49:16]
  assign _T_2574 = ~ _T_2572; // @[LZD.scala 49:27]
  assign _T_2575 = _T_2571 | _T_2574; // @[LZD.scala 49:25]
  assign _T_2576 = _T_2437[3:0]; // @[LZD.scala 49:47]
  assign _T_2577 = _T_2570[3:0]; // @[LZD.scala 49:59]
  assign _T_2578 = _T_2571 ? _T_2576 : _T_2577; // @[LZD.scala 49:35]
  assign _T_2580 = {_T_2573,_T_2575,_T_2578}; // @[Cat.scala 29:58]
  assign _T_2581 = _T_2303[24:0]; // @[LZD.scala 44:32]
  assign _T_2582 = _T_2581[24:9]; // @[LZD.scala 43:32]
  assign _T_2583 = _T_2582[15:8]; // @[LZD.scala 43:32]
  assign _T_2584 = _T_2583[7:4]; // @[LZD.scala 43:32]
  assign _T_2585 = _T_2584[3:2]; // @[LZD.scala 43:32]
  assign _T_2586 = _T_2585 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2587 = _T_2585[1]; // @[LZD.scala 39:21]
  assign _T_2588 = _T_2585[0]; // @[LZD.scala 39:30]
  assign _T_2589 = ~ _T_2588; // @[LZD.scala 39:27]
  assign _T_2590 = _T_2587 | _T_2589; // @[LZD.scala 39:25]
  assign _T_2591 = {_T_2586,_T_2590}; // @[Cat.scala 29:58]
  assign _T_2592 = _T_2584[1:0]; // @[LZD.scala 44:32]
  assign _T_2593 = _T_2592 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2594 = _T_2592[1]; // @[LZD.scala 39:21]
  assign _T_2595 = _T_2592[0]; // @[LZD.scala 39:30]
  assign _T_2596 = ~ _T_2595; // @[LZD.scala 39:27]
  assign _T_2597 = _T_2594 | _T_2596; // @[LZD.scala 39:25]
  assign _T_2598 = {_T_2593,_T_2597}; // @[Cat.scala 29:58]
  assign _T_2599 = _T_2591[1]; // @[Shift.scala 12:21]
  assign _T_2600 = _T_2598[1]; // @[Shift.scala 12:21]
  assign _T_2601 = _T_2599 | _T_2600; // @[LZD.scala 49:16]
  assign _T_2602 = ~ _T_2600; // @[LZD.scala 49:27]
  assign _T_2603 = _T_2599 | _T_2602; // @[LZD.scala 49:25]
  assign _T_2604 = _T_2591[0:0]; // @[LZD.scala 49:47]
  assign _T_2605 = _T_2598[0:0]; // @[LZD.scala 49:59]
  assign _T_2606 = _T_2599 ? _T_2604 : _T_2605; // @[LZD.scala 49:35]
  assign _T_2608 = {_T_2601,_T_2603,_T_2606}; // @[Cat.scala 29:58]
  assign _T_2609 = _T_2583[3:0]; // @[LZD.scala 44:32]
  assign _T_2610 = _T_2609[3:2]; // @[LZD.scala 43:32]
  assign _T_2611 = _T_2610 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2612 = _T_2610[1]; // @[LZD.scala 39:21]
  assign _T_2613 = _T_2610[0]; // @[LZD.scala 39:30]
  assign _T_2614 = ~ _T_2613; // @[LZD.scala 39:27]
  assign _T_2615 = _T_2612 | _T_2614; // @[LZD.scala 39:25]
  assign _T_2616 = {_T_2611,_T_2615}; // @[Cat.scala 29:58]
  assign _T_2617 = _T_2609[1:0]; // @[LZD.scala 44:32]
  assign _T_2618 = _T_2617 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2619 = _T_2617[1]; // @[LZD.scala 39:21]
  assign _T_2620 = _T_2617[0]; // @[LZD.scala 39:30]
  assign _T_2621 = ~ _T_2620; // @[LZD.scala 39:27]
  assign _T_2622 = _T_2619 | _T_2621; // @[LZD.scala 39:25]
  assign _T_2623 = {_T_2618,_T_2622}; // @[Cat.scala 29:58]
  assign _T_2624 = _T_2616[1]; // @[Shift.scala 12:21]
  assign _T_2625 = _T_2623[1]; // @[Shift.scala 12:21]
  assign _T_2626 = _T_2624 | _T_2625; // @[LZD.scala 49:16]
  assign _T_2627 = ~ _T_2625; // @[LZD.scala 49:27]
  assign _T_2628 = _T_2624 | _T_2627; // @[LZD.scala 49:25]
  assign _T_2629 = _T_2616[0:0]; // @[LZD.scala 49:47]
  assign _T_2630 = _T_2623[0:0]; // @[LZD.scala 49:59]
  assign _T_2631 = _T_2624 ? _T_2629 : _T_2630; // @[LZD.scala 49:35]
  assign _T_2633 = {_T_2626,_T_2628,_T_2631}; // @[Cat.scala 29:58]
  assign _T_2634 = _T_2608[2]; // @[Shift.scala 12:21]
  assign _T_2635 = _T_2633[2]; // @[Shift.scala 12:21]
  assign _T_2636 = _T_2634 | _T_2635; // @[LZD.scala 49:16]
  assign _T_2637 = ~ _T_2635; // @[LZD.scala 49:27]
  assign _T_2638 = _T_2634 | _T_2637; // @[LZD.scala 49:25]
  assign _T_2639 = _T_2608[1:0]; // @[LZD.scala 49:47]
  assign _T_2640 = _T_2633[1:0]; // @[LZD.scala 49:59]
  assign _T_2641 = _T_2634 ? _T_2639 : _T_2640; // @[LZD.scala 49:35]
  assign _T_2643 = {_T_2636,_T_2638,_T_2641}; // @[Cat.scala 29:58]
  assign _T_2644 = _T_2582[7:0]; // @[LZD.scala 44:32]
  assign _T_2645 = _T_2644[7:4]; // @[LZD.scala 43:32]
  assign _T_2646 = _T_2645[3:2]; // @[LZD.scala 43:32]
  assign _T_2647 = _T_2646 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2648 = _T_2646[1]; // @[LZD.scala 39:21]
  assign _T_2649 = _T_2646[0]; // @[LZD.scala 39:30]
  assign _T_2650 = ~ _T_2649; // @[LZD.scala 39:27]
  assign _T_2651 = _T_2648 | _T_2650; // @[LZD.scala 39:25]
  assign _T_2652 = {_T_2647,_T_2651}; // @[Cat.scala 29:58]
  assign _T_2653 = _T_2645[1:0]; // @[LZD.scala 44:32]
  assign _T_2654 = _T_2653 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2655 = _T_2653[1]; // @[LZD.scala 39:21]
  assign _T_2656 = _T_2653[0]; // @[LZD.scala 39:30]
  assign _T_2657 = ~ _T_2656; // @[LZD.scala 39:27]
  assign _T_2658 = _T_2655 | _T_2657; // @[LZD.scala 39:25]
  assign _T_2659 = {_T_2654,_T_2658}; // @[Cat.scala 29:58]
  assign _T_2660 = _T_2652[1]; // @[Shift.scala 12:21]
  assign _T_2661 = _T_2659[1]; // @[Shift.scala 12:21]
  assign _T_2662 = _T_2660 | _T_2661; // @[LZD.scala 49:16]
  assign _T_2663 = ~ _T_2661; // @[LZD.scala 49:27]
  assign _T_2664 = _T_2660 | _T_2663; // @[LZD.scala 49:25]
  assign _T_2665 = _T_2652[0:0]; // @[LZD.scala 49:47]
  assign _T_2666 = _T_2659[0:0]; // @[LZD.scala 49:59]
  assign _T_2667 = _T_2660 ? _T_2665 : _T_2666; // @[LZD.scala 49:35]
  assign _T_2669 = {_T_2662,_T_2664,_T_2667}; // @[Cat.scala 29:58]
  assign _T_2670 = _T_2644[3:0]; // @[LZD.scala 44:32]
  assign _T_2671 = _T_2670[3:2]; // @[LZD.scala 43:32]
  assign _T_2672 = _T_2671 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2673 = _T_2671[1]; // @[LZD.scala 39:21]
  assign _T_2674 = _T_2671[0]; // @[LZD.scala 39:30]
  assign _T_2675 = ~ _T_2674; // @[LZD.scala 39:27]
  assign _T_2676 = _T_2673 | _T_2675; // @[LZD.scala 39:25]
  assign _T_2677 = {_T_2672,_T_2676}; // @[Cat.scala 29:58]
  assign _T_2678 = _T_2670[1:0]; // @[LZD.scala 44:32]
  assign _T_2679 = _T_2678 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2680 = _T_2678[1]; // @[LZD.scala 39:21]
  assign _T_2681 = _T_2678[0]; // @[LZD.scala 39:30]
  assign _T_2682 = ~ _T_2681; // @[LZD.scala 39:27]
  assign _T_2683 = _T_2680 | _T_2682; // @[LZD.scala 39:25]
  assign _T_2684 = {_T_2679,_T_2683}; // @[Cat.scala 29:58]
  assign _T_2685 = _T_2677[1]; // @[Shift.scala 12:21]
  assign _T_2686 = _T_2684[1]; // @[Shift.scala 12:21]
  assign _T_2687 = _T_2685 | _T_2686; // @[LZD.scala 49:16]
  assign _T_2688 = ~ _T_2686; // @[LZD.scala 49:27]
  assign _T_2689 = _T_2685 | _T_2688; // @[LZD.scala 49:25]
  assign _T_2690 = _T_2677[0:0]; // @[LZD.scala 49:47]
  assign _T_2691 = _T_2684[0:0]; // @[LZD.scala 49:59]
  assign _T_2692 = _T_2685 ? _T_2690 : _T_2691; // @[LZD.scala 49:35]
  assign _T_2694 = {_T_2687,_T_2689,_T_2692}; // @[Cat.scala 29:58]
  assign _T_2695 = _T_2669[2]; // @[Shift.scala 12:21]
  assign _T_2696 = _T_2694[2]; // @[Shift.scala 12:21]
  assign _T_2697 = _T_2695 | _T_2696; // @[LZD.scala 49:16]
  assign _T_2698 = ~ _T_2696; // @[LZD.scala 49:27]
  assign _T_2699 = _T_2695 | _T_2698; // @[LZD.scala 49:25]
  assign _T_2700 = _T_2669[1:0]; // @[LZD.scala 49:47]
  assign _T_2701 = _T_2694[1:0]; // @[LZD.scala 49:59]
  assign _T_2702 = _T_2695 ? _T_2700 : _T_2701; // @[LZD.scala 49:35]
  assign _T_2704 = {_T_2697,_T_2699,_T_2702}; // @[Cat.scala 29:58]
  assign _T_2705 = _T_2643[3]; // @[Shift.scala 12:21]
  assign _T_2706 = _T_2704[3]; // @[Shift.scala 12:21]
  assign _T_2707 = _T_2705 | _T_2706; // @[LZD.scala 49:16]
  assign _T_2708 = ~ _T_2706; // @[LZD.scala 49:27]
  assign _T_2709 = _T_2705 | _T_2708; // @[LZD.scala 49:25]
  assign _T_2710 = _T_2643[2:0]; // @[LZD.scala 49:47]
  assign _T_2711 = _T_2704[2:0]; // @[LZD.scala 49:59]
  assign _T_2712 = _T_2705 ? _T_2710 : _T_2711; // @[LZD.scala 49:35]
  assign _T_2714 = {_T_2707,_T_2709,_T_2712}; // @[Cat.scala 29:58]
  assign _T_2715 = _T_2581[8:0]; // @[LZD.scala 44:32]
  assign _T_2716 = _T_2715[8:1]; // @[LZD.scala 43:32]
  assign _T_2717 = _T_2716[7:4]; // @[LZD.scala 43:32]
  assign _T_2718 = _T_2717[3:2]; // @[LZD.scala 43:32]
  assign _T_2719 = _T_2718 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2720 = _T_2718[1]; // @[LZD.scala 39:21]
  assign _T_2721 = _T_2718[0]; // @[LZD.scala 39:30]
  assign _T_2722 = ~ _T_2721; // @[LZD.scala 39:27]
  assign _T_2723 = _T_2720 | _T_2722; // @[LZD.scala 39:25]
  assign _T_2724 = {_T_2719,_T_2723}; // @[Cat.scala 29:58]
  assign _T_2725 = _T_2717[1:0]; // @[LZD.scala 44:32]
  assign _T_2726 = _T_2725 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2727 = _T_2725[1]; // @[LZD.scala 39:21]
  assign _T_2728 = _T_2725[0]; // @[LZD.scala 39:30]
  assign _T_2729 = ~ _T_2728; // @[LZD.scala 39:27]
  assign _T_2730 = _T_2727 | _T_2729; // @[LZD.scala 39:25]
  assign _T_2731 = {_T_2726,_T_2730}; // @[Cat.scala 29:58]
  assign _T_2732 = _T_2724[1]; // @[Shift.scala 12:21]
  assign _T_2733 = _T_2731[1]; // @[Shift.scala 12:21]
  assign _T_2734 = _T_2732 | _T_2733; // @[LZD.scala 49:16]
  assign _T_2735 = ~ _T_2733; // @[LZD.scala 49:27]
  assign _T_2736 = _T_2732 | _T_2735; // @[LZD.scala 49:25]
  assign _T_2737 = _T_2724[0:0]; // @[LZD.scala 49:47]
  assign _T_2738 = _T_2731[0:0]; // @[LZD.scala 49:59]
  assign _T_2739 = _T_2732 ? _T_2737 : _T_2738; // @[LZD.scala 49:35]
  assign _T_2741 = {_T_2734,_T_2736,_T_2739}; // @[Cat.scala 29:58]
  assign _T_2742 = _T_2716[3:0]; // @[LZD.scala 44:32]
  assign _T_2743 = _T_2742[3:2]; // @[LZD.scala 43:32]
  assign _T_2744 = _T_2743 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2745 = _T_2743[1]; // @[LZD.scala 39:21]
  assign _T_2746 = _T_2743[0]; // @[LZD.scala 39:30]
  assign _T_2747 = ~ _T_2746; // @[LZD.scala 39:27]
  assign _T_2748 = _T_2745 | _T_2747; // @[LZD.scala 39:25]
  assign _T_2749 = {_T_2744,_T_2748}; // @[Cat.scala 29:58]
  assign _T_2750 = _T_2742[1:0]; // @[LZD.scala 44:32]
  assign _T_2751 = _T_2750 != 2'h0; // @[LZD.scala 39:14]
  assign _T_2752 = _T_2750[1]; // @[LZD.scala 39:21]
  assign _T_2753 = _T_2750[0]; // @[LZD.scala 39:30]
  assign _T_2754 = ~ _T_2753; // @[LZD.scala 39:27]
  assign _T_2755 = _T_2752 | _T_2754; // @[LZD.scala 39:25]
  assign _T_2756 = {_T_2751,_T_2755}; // @[Cat.scala 29:58]
  assign _T_2757 = _T_2749[1]; // @[Shift.scala 12:21]
  assign _T_2758 = _T_2756[1]; // @[Shift.scala 12:21]
  assign _T_2759 = _T_2757 | _T_2758; // @[LZD.scala 49:16]
  assign _T_2760 = ~ _T_2758; // @[LZD.scala 49:27]
  assign _T_2761 = _T_2757 | _T_2760; // @[LZD.scala 49:25]
  assign _T_2762 = _T_2749[0:0]; // @[LZD.scala 49:47]
  assign _T_2763 = _T_2756[0:0]; // @[LZD.scala 49:59]
  assign _T_2764 = _T_2757 ? _T_2762 : _T_2763; // @[LZD.scala 49:35]
  assign _T_2766 = {_T_2759,_T_2761,_T_2764}; // @[Cat.scala 29:58]
  assign _T_2767 = _T_2741[2]; // @[Shift.scala 12:21]
  assign _T_2768 = _T_2766[2]; // @[Shift.scala 12:21]
  assign _T_2769 = _T_2767 | _T_2768; // @[LZD.scala 49:16]
  assign _T_2770 = ~ _T_2768; // @[LZD.scala 49:27]
  assign _T_2771 = _T_2767 | _T_2770; // @[LZD.scala 49:25]
  assign _T_2772 = _T_2741[1:0]; // @[LZD.scala 49:47]
  assign _T_2773 = _T_2766[1:0]; // @[LZD.scala 49:59]
  assign _T_2774 = _T_2767 ? _T_2772 : _T_2773; // @[LZD.scala 49:35]
  assign _T_2776 = {_T_2769,_T_2771,_T_2774}; // @[Cat.scala 29:58]
  assign _T_2777 = _T_2715[0:0]; // @[LZD.scala 44:32]
  assign _T_2779 = _T_2776[3]; // @[Shift.scala 12:21]
  assign _T_2782 = {2'h3,_T_2777}; // @[Cat.scala 29:58]
  assign _T_2783 = _T_2776[2:0]; // @[LZD.scala 55:32]
  assign _T_2784 = _T_2779 ? _T_2783 : _T_2782; // @[LZD.scala 55:20]
  assign _T_2785 = {_T_2779,_T_2784}; // @[Cat.scala 29:58]
  assign _T_2786 = _T_2714[4]; // @[Shift.scala 12:21]
  assign _T_2788 = _T_2714[3:0]; // @[LZD.scala 55:32]
  assign _T_2789 = _T_2786 ? _T_2788 : _T_2785; // @[LZD.scala 55:20]
  assign _T_2790 = {_T_2786,_T_2789}; // @[Cat.scala 29:58]
  assign _T_2791 = _T_2580[5]; // @[Shift.scala 12:21]
  assign _T_2793 = _T_2580[4:0]; // @[LZD.scala 55:32]
  assign _T_2794 = _T_2791 ? _T_2793 : _T_2790; // @[LZD.scala 55:20]
  assign _T_2796 = _T_2302[8]; // @[Shift.scala 12:21]
  assign _T_2799 = {2'h3,_T_2791,_T_2794}; // @[Cat.scala 29:58]
  assign _T_2800 = _T_2302[7:0]; // @[LZD.scala 55:32]
  assign _T_2801 = _T_2796 ? _T_2800 : _T_2799; // @[LZD.scala 55:20]
  assign scaleBias = {1'h1,_T_2796,_T_2801}; // @[Cat.scala 29:58]
  assign _T_2802 = $signed(scaleBias); // @[QuireToPosit.scala 61:53]
  assign _T_2804 = $signed(10'sh11d) + $signed(_T_2802); // @[QuireToPosit.scala 61:41]
  assign realScale = $signed(_T_2804); // @[QuireToPosit.scala 61:41]
  assign underflow = $signed(realScale) < $signed(-10'shf); // @[QuireToPosit.scala 62:41]
  assign overflow = $signed(realScale) > $signed(10'she); // @[QuireToPosit.scala 63:35]
  assign _T_2805 = underflow ? $signed(-10'shf) : $signed(realScale); // @[Mux.scala 87:16]
  assign _T_2806 = overflow ? $signed(10'she) : $signed(_T_2805); // @[Mux.scala 87:16]
  assign _T_2807 = realScale[9:9]; // @[Abs.scala 10:21]
  assign _T_2809 = _T_2807 ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign _T_2810 = $unsigned(realScale); // @[Abs.scala 10:31]
  assign _T_2811 = _T_2809 ^ _T_2810; // @[Abs.scala 10:26]
  assign _GEN_2 = {{9'd0}, _T_2807}; // @[Abs.scala 10:39]
  assign absRealScale = _T_2811 + _GEN_2; // @[Abs.scala 10:39]
  assign _T_2814 = absRealScale < 10'h13a; // @[Shift.scala 16:24]
  assign _T_2815 = absRealScale[8:0]; // @[Shift.scala 17:37]
  assign _T_2816 = _T_2815[8]; // @[Shift.scala 12:21]
  assign _T_2817 = io_quireIn[57:0]; // @[Shift.scala 64:52]
  assign _T_2819 = {_T_2817,256'h0}; // @[Cat.scala 29:58]
  assign _T_2820 = _T_2816 ? _T_2819 : io_quireIn; // @[Shift.scala 64:27]
  assign _T_2821 = _T_2815[7:0]; // @[Shift.scala 66:70]
  assign _T_2822 = _T_2821[7]; // @[Shift.scala 12:21]
  assign _T_2823 = _T_2820[185:0]; // @[Shift.scala 64:52]
  assign _T_2825 = {_T_2823,128'h0}; // @[Cat.scala 29:58]
  assign _T_2826 = _T_2822 ? _T_2825 : _T_2820; // @[Shift.scala 64:27]
  assign _T_2827 = _T_2821[6:0]; // @[Shift.scala 66:70]
  assign _T_2828 = _T_2827[6]; // @[Shift.scala 12:21]
  assign _T_2829 = _T_2826[249:0]; // @[Shift.scala 64:52]
  assign _T_2831 = {_T_2829,64'h0}; // @[Cat.scala 29:58]
  assign _T_2832 = _T_2828 ? _T_2831 : _T_2826; // @[Shift.scala 64:27]
  assign _T_2833 = _T_2827[5:0]; // @[Shift.scala 66:70]
  assign _T_2834 = _T_2833[5]; // @[Shift.scala 12:21]
  assign _T_2835 = _T_2832[281:0]; // @[Shift.scala 64:52]
  assign _T_2837 = {_T_2835,32'h0}; // @[Cat.scala 29:58]
  assign _T_2838 = _T_2834 ? _T_2837 : _T_2832; // @[Shift.scala 64:27]
  assign _T_2839 = _T_2833[4:0]; // @[Shift.scala 66:70]
  assign _T_2840 = _T_2839[4]; // @[Shift.scala 12:21]
  assign _T_2841 = _T_2838[297:0]; // @[Shift.scala 64:52]
  assign _T_2843 = {_T_2841,16'h0}; // @[Cat.scala 29:58]
  assign _T_2844 = _T_2840 ? _T_2843 : _T_2838; // @[Shift.scala 64:27]
  assign _T_2845 = _T_2839[3:0]; // @[Shift.scala 66:70]
  assign _T_2846 = _T_2845[3]; // @[Shift.scala 12:21]
  assign _T_2847 = _T_2844[305:0]; // @[Shift.scala 64:52]
  assign _T_2849 = {_T_2847,8'h0}; // @[Cat.scala 29:58]
  assign _T_2850 = _T_2846 ? _T_2849 : _T_2844; // @[Shift.scala 64:27]
  assign _T_2851 = _T_2845[2:0]; // @[Shift.scala 66:70]
  assign _T_2852 = _T_2851[2]; // @[Shift.scala 12:21]
  assign _T_2853 = _T_2850[309:0]; // @[Shift.scala 64:52]
  assign _T_2855 = {_T_2853,4'h0}; // @[Cat.scala 29:58]
  assign _T_2856 = _T_2852 ? _T_2855 : _T_2850; // @[Shift.scala 64:27]
  assign _T_2857 = _T_2851[1:0]; // @[Shift.scala 66:70]
  assign _T_2858 = _T_2857[1]; // @[Shift.scala 12:21]
  assign _T_2859 = _T_2856[311:0]; // @[Shift.scala 64:52]
  assign _T_2861 = {_T_2859,2'h0}; // @[Cat.scala 29:58]
  assign _T_2862 = _T_2858 ? _T_2861 : _T_2856; // @[Shift.scala 64:27]
  assign _T_2863 = _T_2857[0:0]; // @[Shift.scala 66:70]
  assign _T_2865 = _T_2862[312:0]; // @[Shift.scala 64:52]
  assign _T_2866 = {_T_2865,1'h0}; // @[Cat.scala 29:58]
  assign _T_2867 = _T_2863 ? _T_2866 : _T_2862; // @[Shift.scala 64:27]
  assign quireLeftShift = _T_2814 ? _T_2867 : 314'h0; // @[Shift.scala 16:10]
  assign _T_2872 = io_quireIn[313:256]; // @[Shift.scala 77:66]
  assign _T_2873 = {256'h0,_T_2872}; // @[Cat.scala 29:58]
  assign _T_2874 = _T_2816 ? _T_2873 : io_quireIn; // @[Shift.scala 77:22]
  assign _T_2878 = _T_2874[313:128]; // @[Shift.scala 77:66]
  assign _T_2879 = {128'h0,_T_2878}; // @[Cat.scala 29:58]
  assign _T_2880 = _T_2822 ? _T_2879 : _T_2874; // @[Shift.scala 77:22]
  assign _T_2884 = _T_2880[313:64]; // @[Shift.scala 77:66]
  assign _T_2885 = {64'h0,_T_2884}; // @[Cat.scala 29:58]
  assign _T_2886 = _T_2828 ? _T_2885 : _T_2880; // @[Shift.scala 77:22]
  assign _T_2890 = _T_2886[313:32]; // @[Shift.scala 77:66]
  assign _T_2891 = {32'h0,_T_2890}; // @[Cat.scala 29:58]
  assign _T_2892 = _T_2834 ? _T_2891 : _T_2886; // @[Shift.scala 77:22]
  assign _T_2896 = _T_2892[313:16]; // @[Shift.scala 77:66]
  assign _T_2897 = {16'h0,_T_2896}; // @[Cat.scala 29:58]
  assign _T_2898 = _T_2840 ? _T_2897 : _T_2892; // @[Shift.scala 77:22]
  assign _T_2902 = _T_2898[313:8]; // @[Shift.scala 77:66]
  assign _T_2903 = {8'h0,_T_2902}; // @[Cat.scala 29:58]
  assign _T_2904 = _T_2846 ? _T_2903 : _T_2898; // @[Shift.scala 77:22]
  assign _T_2908 = _T_2904[313:4]; // @[Shift.scala 77:66]
  assign _T_2909 = {4'h0,_T_2908}; // @[Cat.scala 29:58]
  assign _T_2910 = _T_2852 ? _T_2909 : _T_2904; // @[Shift.scala 77:22]
  assign _T_2914 = _T_2910[313:2]; // @[Shift.scala 77:66]
  assign _T_2915 = {2'h0,_T_2914}; // @[Cat.scala 29:58]
  assign _T_2916 = _T_2858 ? _T_2915 : _T_2910; // @[Shift.scala 77:22]
  assign _T_2919 = _T_2916[313:1]; // @[Shift.scala 77:66]
  assign _T_2920 = {1'h0,_T_2919}; // @[Cat.scala 29:58]
  assign _T_2921 = _T_2863 ? _T_2920 : _T_2916; // @[Shift.scala 77:22]
  assign quireRightShift = _T_2814 ? _T_2921 : 314'h0; // @[Shift.scala 27:10]
  assign _T_2923 = quireLeftShift[27:13]; // @[QuireToPosit.scala 89:49]
  assign _T_2924 = quireLeftShift[12:0]; // @[QuireToPosit.scala 90:127]
  assign _T_2925 = _T_2924 != 13'h0; // @[QuireToPosit.scala 90:154]
  assign realFGRSTmp1 = {_T_2923,_T_2925}; // @[Cat.scala 29:58]
  assign _T_2926 = quireRightShift[27:13]; // @[QuireToPosit.scala 91:50]
  assign _T_2927 = quireRightShift[12:0]; // @[QuireToPosit.scala 92:128]
  assign _T_2928 = _T_2927 != 13'h0; // @[QuireToPosit.scala 92:155]
  assign realFGRSTmp2 = {_T_2926,_T_2928}; // @[Cat.scala 29:58]
  assign realFGRS = _T_2807 ? realFGRSTmp1 : realFGRSTmp2; // @[QuireToPosit.scala 93:34]
  assign outRawFloat_fraction = realFGRS[15:3]; // @[QuireToPosit.scala 95:46]
  assign outRawFloat_grs = realFGRS[2:0]; // @[QuireToPosit.scala 96:46]
  assign _GEN_3 = _T_2806[4:0]; // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  assign outRawFloat_scale = $signed(_GEN_3); // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  assign _T_2934 = outRawFloat_scale[4:4]; // @[convert.scala 49:36]
  assign _T_2936 = ~ outRawFloat_scale; // @[convert.scala 50:36]
  assign _T_2937 = $signed(_T_2936); // @[convert.scala 50:36]
  assign _T_2938 = _T_2934 ? $signed(_T_2937) : $signed(outRawFloat_scale); // @[convert.scala 50:28]
  assign _T_2939 = _T_2934 ^ _T_2; // @[convert.scala 51:31]
  assign _T_2940 = ~ _T_2939; // @[convert.scala 53:34]
  assign _T_2943 = {_T_2940,_T_2939,outRawFloat_fraction,outRawFloat_grs}; // @[Cat.scala 29:58]
  assign _T_2944 = $unsigned(_T_2938); // @[Shift.scala 39:17]
  assign _T_2945 = _T_2944 < 5'h12; // @[Shift.scala 39:24]
  assign _T_2947 = _T_2943[17:16]; // @[Shift.scala 90:30]
  assign _T_2948 = _T_2943[15:0]; // @[Shift.scala 90:48]
  assign _T_2949 = _T_2948 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_4 = {{1'd0}, _T_2949}; // @[Shift.scala 90:39]
  assign _T_2950 = _T_2947 | _GEN_4; // @[Shift.scala 90:39]
  assign _T_2951 = _T_2944[4]; // @[Shift.scala 12:21]
  assign _T_2952 = _T_2943[17]; // @[Shift.scala 12:21]
  assign _T_2954 = _T_2952 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_2955 = {_T_2954,_T_2950}; // @[Cat.scala 29:58]
  assign _T_2956 = _T_2951 ? _T_2955 : _T_2943; // @[Shift.scala 91:22]
  assign _T_2957 = _T_2944[3:0]; // @[Shift.scala 92:77]
  assign _T_2958 = _T_2956[17:8]; // @[Shift.scala 90:30]
  assign _T_2959 = _T_2956[7:0]; // @[Shift.scala 90:48]
  assign _T_2960 = _T_2959 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_5 = {{9'd0}, _T_2960}; // @[Shift.scala 90:39]
  assign _T_2961 = _T_2958 | _GEN_5; // @[Shift.scala 90:39]
  assign _T_2962 = _T_2957[3]; // @[Shift.scala 12:21]
  assign _T_2963 = _T_2956[17]; // @[Shift.scala 12:21]
  assign _T_2965 = _T_2963 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_2966 = {_T_2965,_T_2961}; // @[Cat.scala 29:58]
  assign _T_2967 = _T_2962 ? _T_2966 : _T_2956; // @[Shift.scala 91:22]
  assign _T_2968 = _T_2957[2:0]; // @[Shift.scala 92:77]
  assign _T_2969 = _T_2967[17:4]; // @[Shift.scala 90:30]
  assign _T_2970 = _T_2967[3:0]; // @[Shift.scala 90:48]
  assign _T_2971 = _T_2970 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_6 = {{13'd0}, _T_2971}; // @[Shift.scala 90:39]
  assign _T_2972 = _T_2969 | _GEN_6; // @[Shift.scala 90:39]
  assign _T_2973 = _T_2968[2]; // @[Shift.scala 12:21]
  assign _T_2974 = _T_2967[17]; // @[Shift.scala 12:21]
  assign _T_2976 = _T_2974 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_2977 = {_T_2976,_T_2972}; // @[Cat.scala 29:58]
  assign _T_2978 = _T_2973 ? _T_2977 : _T_2967; // @[Shift.scala 91:22]
  assign _T_2979 = _T_2968[1:0]; // @[Shift.scala 92:77]
  assign _T_2980 = _T_2978[17:2]; // @[Shift.scala 90:30]
  assign _T_2981 = _T_2978[1:0]; // @[Shift.scala 90:48]
  assign _T_2982 = _T_2981 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_7 = {{15'd0}, _T_2982}; // @[Shift.scala 90:39]
  assign _T_2983 = _T_2980 | _GEN_7; // @[Shift.scala 90:39]
  assign _T_2984 = _T_2979[1]; // @[Shift.scala 12:21]
  assign _T_2985 = _T_2978[17]; // @[Shift.scala 12:21]
  assign _T_2987 = _T_2985 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_2988 = {_T_2987,_T_2983}; // @[Cat.scala 29:58]
  assign _T_2989 = _T_2984 ? _T_2988 : _T_2978; // @[Shift.scala 91:22]
  assign _T_2990 = _T_2979[0:0]; // @[Shift.scala 92:77]
  assign _T_2991 = _T_2989[17:1]; // @[Shift.scala 90:30]
  assign _T_2992 = _T_2989[0:0]; // @[Shift.scala 90:48]
  assign _GEN_8 = {{16'd0}, _T_2992}; // @[Shift.scala 90:39]
  assign _T_2994 = _T_2991 | _GEN_8; // @[Shift.scala 90:39]
  assign _T_2996 = _T_2989[17]; // @[Shift.scala 12:21]
  assign _T_2997 = {_T_2996,_T_2994}; // @[Cat.scala 29:58]
  assign _T_2998 = _T_2990 ? _T_2997 : _T_2989; // @[Shift.scala 91:22]
  assign _T_3001 = _T_2952 ? 18'h3ffff : 18'h0; // @[Bitwise.scala 71:12]
  assign _T_3002 = _T_2945 ? _T_2998 : _T_3001; // @[Shift.scala 39:10]
  assign _T_3003 = _T_3002[3]; // @[convert.scala 55:31]
  assign _T_3004 = _T_3002[2]; // @[convert.scala 56:31]
  assign _T_3005 = _T_3002[1]; // @[convert.scala 57:31]
  assign _T_3006 = _T_3002[0]; // @[convert.scala 58:31]
  assign _T_3007 = _T_3002[17:3]; // @[convert.scala 59:69]
  assign _T_3008 = _T_3007 != 15'h0; // @[convert.scala 59:81]
  assign _T_3009 = ~ _T_3008; // @[convert.scala 59:50]
  assign _T_3011 = _T_3007 == 15'h7fff; // @[convert.scala 60:81]
  assign _T_3012 = _T_3003 | _T_3005; // @[convert.scala 61:44]
  assign _T_3013 = _T_3012 | _T_3006; // @[convert.scala 61:52]
  assign _T_3014 = _T_3004 & _T_3013; // @[convert.scala 61:36]
  assign _T_3015 = ~ _T_3011; // @[convert.scala 62:63]
  assign _T_3016 = _T_3015 & _T_3014; // @[convert.scala 62:103]
  assign _T_3017 = _T_3009 | _T_3016; // @[convert.scala 62:60]
  assign _GEN_9 = {{14'd0}, _T_3017}; // @[convert.scala 63:56]
  assign _T_3020 = _T_3007 + _GEN_9; // @[convert.scala 63:56]
  assign _T_3021 = {_T_2,_T_3020}; // @[Cat.scala 29:58]
  assign io_positOut = _T_3029; // @[QuireToPosit.scala 101:15]
  assign io_outValid = _T_3025; // @[QuireToPosit.scala 100:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_3025 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_3029 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_3025 <= 1'h0;
    end else begin
      _T_3025 <= io_inValid;
    end
    if (io_inValid) begin
      if (outRawFloat_isNaR) begin
        _T_3029 <= 16'h8000;
      end else begin
        if (outRawFloat_isZero) begin
          _T_3029 <= 16'h0;
        end else begin
          _T_3029 <= _T_3021;
        end
      end
    end
  end
endmodule
